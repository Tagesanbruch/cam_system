// Verilog netlist created by Tang Dynasty v6.0.122666
// Wed Oct 16 22:27:55 2024

`timescale 1ns / 1ps
module AnlCORDIC_sqrt
  (
  clk,
  num,
  rst,
  start,
  done,
  sqrt
  );

  input clk;
  input [20:0] num;
  input rst;
  input start;
  output done;
  output [20:0] sqrt;

  parameter COMPENSATION = "No Compensation";
  parameter ITERATION = 10;
  parameter PRECISION = 20;
  parameter SCALED = 0;
  // localparam W_CNT = 4;
  // localparam W_SFT = 5;
  wire [20:0] al_92abc73b;
  wire [20:0] al_5a529b34;
  wire [20:0] al_6d90eb23;
  wire [3:0] al_b029b709;
  wire [20:0] al_c21a53a9;
  wire  al_b2a2e5ce;
  wire  al_fe92b9c9;
  wire  al_14573418;
  wire  al_1f8ac62a;
  wire  al_1e89e993;
  wire  al_b81bed99;
  wire  al_64d5f40e;
  wire  al_fb75ed64;
  wire  al_81b0c7fb;
  wire  al_f33a944d;
  wire  al_a65c875a;
  wire  al_da2dd23a;
  wire  al_86dcc04b;
  wire  al_43cf9c51;
  wire  al_312b9047;
  wire  al_6bd399c8;
  wire  al_7406b7f;
  wire  al_68be76e6;
  wire  al_f3ac4ff4;
  wire  al_462198a;
  wire  al_2ec9e601;
  wire  al_c9156751;
  wire  al_ded0a164;
  wire  al_c6dd6de;
  wire  al_db11fb22;
  wire  al_3f457ae0;
  wire  al_8f7d8418;
  wire  al_c4b36f25;
  wire  al_a6f911fa;
  wire  al_3a11d010;
  wire  al_5976b207;
  wire  al_1aa4ae3e;
  wire  al_da6a2c78;
  wire  al_124b3a01;
  wire  al_f35b497d;
  wire  al_7f73cd24;
  wire  al_da90d6e3;
  wire  al_b1cdfbfa;
  wire  al_695678a9;
  wire  al_9be05a01;
  wire  al_cbac66be;
  wire  al_4b0ede28;
  wire  al_24ebd63f;
  wire  al_8a0179a4;
  wire  al_d7a13544;
  wire  al_a4ba3987;
  wire  al_b6c514a3;
  wire  al_4559aa8f;
  wire  al_60425dcb;
  wire  al_dacf88bd;
  wire  al_a614d965;
  wire  al_54282d1f;
  wire  al_a6672972;
  wire  al_15a841b9;
  wire  al_3dc3e1bb;
  wire  al_76d214f0;
  wire  al_fdf9855e;
  wire  al_83c825e4;
  wire  al_babeab3;
  wire  al_a67e0f03;
  wire  al_ab2fd291;
  wire  al_a60487f4;
  wire  al_dd9cb274;
  wire  al_f0c918f2;
  wire  al_b050724b;
  wire  al_f3539fe0;
  wire [4:0] al_e01c36e7;
  wire [4:0] al_338a517;
  wire [20:0] al_6de4c23f;
  wire [22:0] al_16357ce4;
  wire [22:0] al_f8bbbf13;
  wire [19:0] al_378a1ee4;
  wire [22:0] al_8ff04cfd;
  wire [22:0] al_d65643ad;
  wire [22:0] al_7b2fe207;
  wire [22:0] al_da03ca6b;
  wire [22:0] al_cbee0ff9;
  wire [22:0] al_de90ce1b;
  wire [22:0] al_c968c273;
  wire [22:0] al_19b5d2a2;
  wire al_fcc7c8eb;
  wire al_bfc62871;
  wire al_a83efe58;
  wire al_9c438f85;
  wire al_6e4658ce;
  wire al_d13cd7d5;
  wire al_a7c1a5ec;
  wire al_904f176;
  wire al_ae05c008;
  wire al_583c41b;
  wire al_56a70e01;
  wire al_a5de408f;
  wire al_2231b599;
  wire al_78a16a1;
  wire al_5c2d1b17;
  wire al_c90b7a29;
  wire al_c875ca4a;
  wire al_fc7719ff;
  wire al_36250f57;
  wire al_a5eacf43;
  wire al_7534d24c;
  wire al_1f0013fa;
  wire al_99f44ac;
  wire al_d0045161;
  wire al_16c52ec8;
  wire al_af21225a;
  wire al_8ba9d093;
  wire al_d2041f17;
  wire al_477219c8;
  wire al_df76032a;
  wire al_ff46c763;
  wire al_b24dfd83;
  wire al_c118201a;
  wire al_d6beb4eb;
  wire al_49771648;
  wire al_ebd6c8eb;
  wire al_4504bc33;
  wire al_3b7fed09;
  wire al_545f7ecb;
  wire al_26f5ffe0;
  wire al_c7cb74b5;
  wire al_61d1252c;
  wire al_bb682414;
  wire al_a5340e3c;
  wire al_a3421794;
  wire al_74db697d;
  wire al_5415e4e8;
  wire al_3b78300a;
  wire al_cfbcfa66;
  wire al_32aef229;
  wire al_ef2c5c41;
  wire al_74a93460;
  wire al_44bf9465;
  wire al_b9f06911;
  wire al_dbc76591;
  wire al_90ab3623;
  wire al_58a71ac4;
  wire al_bcd67f57;
  wire al_d7d54632;
  wire al_16ac7bbd;
  wire al_b1b6696e;
  wire al_3f0678ce;
  wire al_848f0c09;
  wire al_ad6322d2;
  wire al_d2549e3b;
  wire al_a47b1084;
  wire al_2dff9c9f;
  wire al_82338500;
  wire al_5669eee7;
  wire al_653faf9;
  wire al_337720e7;
  wire al_e013aab4;
  wire al_304d439a;
  wire al_7adb5007;
  wire al_d5ae2d7f;
  wire al_6c0808;
  wire al_ae0a6293;
  wire al_d07a623a;
  wire al_126bbf82;
  wire al_1aac3445;
  wire al_f5516224;
  wire al_91108e0e;
  wire al_a4e1781b;
  wire al_dc44be48;
  wire al_d8dd00e3;
  wire al_a0bad8f5;
  wire al_c93e73fa;
  wire al_6ea85cef;
  wire al_52616de9;
  wire al_ec1119c9;
  wire al_77f3553d;
  wire al_6299424f;
  wire al_ea5880d3;
  wire al_bbe9aae2;
  wire al_d9ef6091;
  wire al_7109a3cd;
  wire al_f1bac0a6;
  wire al_61c118b2;
  wire al_9bb03b7;
  wire al_d6d4ff9e;
  wire al_b6ba68ca;
  wire al_3c3af6b1;
  wire al_c7e7c580;
  wire al_a93520ae;
  wire al_81c04c9c;
  wire al_f584a17a;
  wire al_5d663e44;
  wire al_27011e73;
  wire al_4c0f5956;
  wire al_e0589574;
  wire al_12f8fb3c;
  wire al_3c4a6475;
  wire al_9fa575eb;
  wire al_d3327d96;
  wire al_412f61d0;
  wire al_3b62f46f;
  wire al_5d141531;
  wire al_67aa9deb;
  wire al_3697e743;
  wire al_3d62c9fe;
  wire al_81a11f5a;
  wire al_461d7931;
  wire al_42fa3115;
  wire al_e2e350ce;
  wire al_a4c5989a;
  wire al_c34f1a86;
  wire al_11b32505;
  wire al_2a2e2537;
  wire al_b4044579;
  wire al_4090ecdb;
  wire al_b1c2c144;
  wire al_60d662e6;
  wire al_687e23a0;
  wire al_b5c4be4e;
  wire al_f1e4a7a7;
  wire al_e2931770;
  wire al_4821ff7f;
  wire al_712165e6;
  wire al_1749b8de;
  wire al_593536de;
  wire al_8f6c5547;
  wire al_ff178429;
  wire al_a46cb2d7;
  wire al_4e7e9688;
  wire al_f7b167;
  wire al_9ea00fd2;
  wire al_a7063677;
  wire al_fa2e23e1;
  wire al_91a73912;
  wire al_e1b97ac;
  wire al_8b1fe6d5;
  wire al_2b66b96f;
  wire al_6067595f;
  wire al_75977872;
  wire al_d3758072;
  wire al_6b3505b5;
  wire al_fa86226a;
  wire al_500d0cf0;
  wire al_8563d1ec;
  wire al_3123bab1;
  wire al_a67b2030;
  wire al_a980305;
  wire al_c3ad1f75;
  wire al_788d5b83;
  wire al_ae3fe1e5;
  wire al_1823807d;
  wire al_36c58aac;
  wire al_45db9cb5;
  wire al_4fb683a3;
  wire al_8c06569d;
  wire al_5c9f255f;
  wire al_696d4179;
  wire al_6979d612;
  wire al_8bf09624;
  wire al_db63ae90;
  wire al_57322515;
  wire al_e75a278b;
  wire al_3261239f;
  wire al_a2611309;
  wire al_3896e32f;
  wire al_1ea08bcc;
  wire al_534eeb32;
  wire al_66f5623c;
  wire al_f5e8ffb7;
  wire al_de41ded2;
  wire al_803879c7;
  wire al_6f8464f;
  wire al_3127e1e8;
  wire al_c162c2a5;

  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_6df20a54 (
    .a(1'b0),
    .o({al_fcc7c8eb,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8d80c396 (
    .a(al_92abc73b[1]),
    .b(1'b1),
    .c(al_fcc7c8eb),
    .o({al_bfc62871,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_22dfbf6 (
    .a(al_92abc73b[2]),
    .b(1'b0),
    .c(al_bfc62871),
    .o({al_a83efe58,al_378a1ee4[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b6ce109b (
    .a(al_92abc73b[3]),
    .b(1'b1),
    .c(al_a83efe58),
    .o({al_9c438f85,al_378a1ee4[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3be7cdd2 (
    .a(al_92abc73b[4]),
    .b(1'b0),
    .c(al_9c438f85),
    .o({al_6e4658ce,al_378a1ee4[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_abc5c8fc (
    .a(al_92abc73b[5]),
    .b(1'b0),
    .c(al_6e4658ce),
    .o({al_d13cd7d5,al_378a1ee4[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_35dee330 (
    .a(al_92abc73b[6]),
    .b(1'b0),
    .c(al_d13cd7d5),
    .o({al_a7c1a5ec,al_378a1ee4[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a6a3e0a0 (
    .a(al_92abc73b[7]),
    .b(1'b0),
    .c(al_a7c1a5ec),
    .o({al_904f176,al_378a1ee4[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cea749b0 (
    .a(al_92abc73b[8]),
    .b(1'b1),
    .c(al_904f176),
    .o({al_ae05c008,al_378a1ee4[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6d66ee19 (
    .a(al_92abc73b[9]),
    .b(1'b0),
    .c(al_ae05c008),
    .o({al_583c41b,al_378a1ee4[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3bbe2c91 (
    .a(al_92abc73b[10]),
    .b(1'b1),
    .c(al_583c41b),
    .o({al_56a70e01,al_378a1ee4[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_41d36f2b (
    .a(al_92abc73b[11]),
    .b(1'b0),
    .c(al_56a70e01),
    .o({al_a5de408f,al_378a1ee4[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8b54afaf (
    .a(al_92abc73b[12]),
    .b(1'b1),
    .c(al_a5de408f),
    .o({al_2231b599,al_378a1ee4[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_90b1a19d (
    .a(al_92abc73b[13]),
    .b(1'b0),
    .c(al_2231b599),
    .o({al_78a16a1,al_378a1ee4[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e56607bb (
    .a(al_92abc73b[14]),
    .b(1'b1),
    .c(al_78a16a1),
    .o({al_5c2d1b17,al_378a1ee4[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4e97fc42 (
    .a(al_92abc73b[15]),
    .b(1'b1),
    .c(al_5c2d1b17),
    .o({al_c90b7a29,al_378a1ee4[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_29d0fe45 (
    .a(al_92abc73b[16]),
    .b(1'b1),
    .c(al_c90b7a29),
    .o({al_c875ca4a,al_378a1ee4[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f04e2943 (
    .a(al_92abc73b[17]),
    .b(1'b0),
    .c(al_c875ca4a),
    .o({al_fc7719ff,al_378a1ee4[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4566af8 (
    .a(al_92abc73b[18]),
    .b(1'b1),
    .c(al_fc7719ff),
    .o({al_36250f57,al_378a1ee4[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_33f9013e (
    .a(al_92abc73b[19]),
    .b(1'b0),
    .c(al_36250f57),
    .o({al_a5eacf43,al_378a1ee4[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4c65cb8e (
    .a(al_92abc73b[20]),
    .b(1'b0),
    .c(al_a5eacf43),
    .o({al_7534d24c,al_378a1ee4[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_da4d991f (
    .c(al_7534d24c),
    .o({open_n6,al_6f8464f}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c22ee456 (
    .a(al_16357ce4[7]),
    .b(al_19b5d2a2[7]),
    .c(al_477219c8),
    .o({al_df76032a,al_d65643ad[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d4f8c6b2 (
    .a(al_16357ce4[8]),
    .b(al_19b5d2a2[8]),
    .c(al_df76032a),
    .o({al_ff46c763,al_d65643ad[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_251c9501 (
    .a(al_16357ce4[9]),
    .b(al_19b5d2a2[9]),
    .c(al_ff46c763),
    .o({al_b24dfd83,al_d65643ad[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b10f851 (
    .a(al_16357ce4[10]),
    .b(al_19b5d2a2[10]),
    .c(al_b24dfd83),
    .o({al_c118201a,al_d65643ad[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f6074d25 (
    .a(al_16357ce4[11]),
    .b(al_19b5d2a2[11]),
    .c(al_c118201a),
    .o({al_d6beb4eb,al_d65643ad[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fa8db078 (
    .a(al_16357ce4[12]),
    .b(al_19b5d2a2[12]),
    .c(al_d6beb4eb),
    .o({al_49771648,al_d65643ad[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_77855a53 (
    .a(al_16357ce4[13]),
    .b(al_19b5d2a2[13]),
    .c(al_49771648),
    .o({al_ebd6c8eb,al_d65643ad[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e3fa0367 (
    .a(al_16357ce4[14]),
    .b(al_19b5d2a2[14]),
    .c(al_ebd6c8eb),
    .o({al_4504bc33,al_d65643ad[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f953a96c (
    .a(al_16357ce4[15]),
    .b(al_19b5d2a2[15]),
    .c(al_4504bc33),
    .o({al_3b7fed09,al_d65643ad[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_65c8a090 (
    .a(al_16357ce4[16]),
    .b(al_19b5d2a2[16]),
    .c(al_3b7fed09),
    .o({al_545f7ecb,al_d65643ad[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_542d5c78 (
    .a(1'b0),
    .o({al_1f0013fa,open_n9}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_53b7c044 (
    .a(al_16357ce4[17]),
    .b(al_19b5d2a2[17]),
    .c(al_545f7ecb),
    .o({al_26f5ffe0,al_d65643ad[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d4fabdf4 (
    .a(al_16357ce4[18]),
    .b(al_19b5d2a2[18]),
    .c(al_26f5ffe0),
    .o({al_c7cb74b5,al_d65643ad[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4c333d3d (
    .a(al_16357ce4[19]),
    .b(al_19b5d2a2[19]),
    .c(al_c7cb74b5),
    .o({al_61d1252c,al_d65643ad[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ad500350 (
    .a(al_16357ce4[20]),
    .b(al_19b5d2a2[20]),
    .c(al_61d1252c),
    .o({al_bb682414,al_d65643ad[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d576b9a4 (
    .a(al_16357ce4[21]),
    .b(al_19b5d2a2[21]),
    .c(al_bb682414),
    .o({al_a5340e3c,al_d65643ad[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e0e9c2f2 (
    .a(al_16357ce4[22]),
    .b(al_19b5d2a2[21]),
    .c(al_a5340e3c),
    .o({open_n10,al_d65643ad[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a685a1be (
    .a(al_16357ce4[0]),
    .b(al_19b5d2a2[0]),
    .c(al_1f0013fa),
    .o({al_99f44ac,al_d65643ad[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cda14380 (
    .a(al_16357ce4[1]),
    .b(al_19b5d2a2[1]),
    .c(al_99f44ac),
    .o({al_d0045161,al_d65643ad[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f54c3dbb (
    .a(al_16357ce4[2]),
    .b(al_19b5d2a2[2]),
    .c(al_d0045161),
    .o({al_16c52ec8,al_d65643ad[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c9b145c3 (
    .a(al_16357ce4[3]),
    .b(al_19b5d2a2[3]),
    .c(al_16c52ec8),
    .o({al_af21225a,al_d65643ad[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_85743617 (
    .a(al_16357ce4[4]),
    .b(al_19b5d2a2[4]),
    .c(al_af21225a),
    .o({al_8ba9d093,al_d65643ad[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ad670f93 (
    .a(al_16357ce4[5]),
    .b(al_19b5d2a2[5]),
    .c(al_8ba9d093),
    .o({al_d2041f17,al_d65643ad[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ec16458c (
    .a(al_16357ce4[6]),
    .b(al_19b5d2a2[6]),
    .c(al_d2041f17),
    .o({al_477219c8,al_d65643ad[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5a77c71d (
    .a(al_da03ca6b[7]),
    .b(al_7b2fe207[7]),
    .c(al_74a93460),
    .o({al_44bf9465,al_c968c273[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6113318c (
    .a(al_da03ca6b[8]),
    .b(al_7b2fe207[8]),
    .c(al_44bf9465),
    .o({al_b9f06911,al_c968c273[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1ba0daa2 (
    .a(al_da03ca6b[9]),
    .b(al_7b2fe207[9]),
    .c(al_b9f06911),
    .o({al_dbc76591,al_c968c273[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4ff26d7e (
    .a(al_da03ca6b[10]),
    .b(al_7b2fe207[10]),
    .c(al_dbc76591),
    .o({al_90ab3623,al_c968c273[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b257243f (
    .a(al_da03ca6b[11]),
    .b(al_7b2fe207[11]),
    .c(al_90ab3623),
    .o({al_58a71ac4,al_c968c273[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ce1cc971 (
    .a(al_da03ca6b[12]),
    .b(al_7b2fe207[12]),
    .c(al_58a71ac4),
    .o({al_bcd67f57,al_c968c273[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e3dc02b8 (
    .a(al_da03ca6b[13]),
    .b(al_7b2fe207[13]),
    .c(al_bcd67f57),
    .o({al_d7d54632,al_c968c273[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9fa2507d (
    .a(al_da03ca6b[14]),
    .b(al_7b2fe207[14]),
    .c(al_d7d54632),
    .o({al_16ac7bbd,al_c968c273[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f7236576 (
    .a(al_da03ca6b[15]),
    .b(al_7b2fe207[15]),
    .c(al_16ac7bbd),
    .o({al_b1b6696e,al_c968c273[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d5b75486 (
    .a(al_da03ca6b[16]),
    .b(al_7b2fe207[16]),
    .c(al_b1b6696e),
    .o({al_3f0678ce,al_c968c273[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_61c46b5d (
    .a(1'b0),
    .o({al_a3421794,open_n13}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2785c3f1 (
    .a(al_da03ca6b[17]),
    .b(al_7b2fe207[17]),
    .c(al_3f0678ce),
    .o({al_848f0c09,al_c968c273[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cb06c7bc (
    .a(al_da03ca6b[18]),
    .b(al_7b2fe207[18]),
    .c(al_848f0c09),
    .o({al_ad6322d2,al_c968c273[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ec350d83 (
    .a(al_da03ca6b[19]),
    .b(al_7b2fe207[19]),
    .c(al_ad6322d2),
    .o({al_d2549e3b,al_c968c273[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c2dfa21e (
    .a(al_da03ca6b[20]),
    .b(al_7b2fe207[20]),
    .c(al_d2549e3b),
    .o({al_a47b1084,al_c968c273[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_19307c7a (
    .a(al_da03ca6b[21]),
    .b(al_7b2fe207[21]),
    .c(al_a47b1084),
    .o({al_2dff9c9f,al_c968c273[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cae2bf94 (
    .a(al_da03ca6b[22]),
    .b(al_7b2fe207[21]),
    .c(al_2dff9c9f),
    .o({open_n14,al_c968c273[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9c5c9996 (
    .a(al_da03ca6b[0]),
    .b(al_7b2fe207[0]),
    .c(al_a3421794),
    .o({al_74db697d,al_c968c273[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c04cf982 (
    .a(al_da03ca6b[1]),
    .b(al_7b2fe207[1]),
    .c(al_74db697d),
    .o({al_5415e4e8,al_c968c273[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f1d55d58 (
    .a(al_da03ca6b[2]),
    .b(al_7b2fe207[2]),
    .c(al_5415e4e8),
    .o({al_3b78300a,al_c968c273[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_212b0a99 (
    .a(al_da03ca6b[3]),
    .b(al_7b2fe207[3]),
    .c(al_3b78300a),
    .o({al_cfbcfa66,al_c968c273[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4a0be642 (
    .a(al_da03ca6b[4]),
    .b(al_7b2fe207[4]),
    .c(al_cfbcfa66),
    .o({al_32aef229,al_c968c273[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9d22fee2 (
    .a(al_da03ca6b[5]),
    .b(al_7b2fe207[5]),
    .c(al_32aef229),
    .o({al_ef2c5c41,al_c968c273[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a9fc3313 (
    .a(al_da03ca6b[6]),
    .b(al_7b2fe207[6]),
    .c(al_ef2c5c41),
    .o({al_74a93460,al_c968c273[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_bcb73af7 (
    .a(1'b0),
    .o({al_e2e350ce,open_n17}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17fb46fe (
    .a(al_92abc73b[1]),
    .b(1'b1),
    .c(al_e2e350ce),
    .o({al_a4c5989a,open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_84c18b6d (
    .a(al_92abc73b[2]),
    .b(1'b0),
    .c(al_a4c5989a),
    .o({al_c34f1a86,open_n19}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dd32fe7c (
    .a(al_92abc73b[3]),
    .b(1'b1),
    .c(al_c34f1a86),
    .o({al_11b32505,al_5a529b34[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d535d783 (
    .a(al_92abc73b[4]),
    .b(1'b0),
    .c(al_11b32505),
    .o({al_2a2e2537,al_5a529b34[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_47e8f6cc (
    .a(al_92abc73b[5]),
    .b(1'b0),
    .c(al_2a2e2537),
    .o({al_b4044579,al_5a529b34[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d8de1e47 (
    .a(al_92abc73b[6]),
    .b(1'b0),
    .c(al_b4044579),
    .o({al_4090ecdb,al_5a529b34[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_70762dc4 (
    .a(al_92abc73b[7]),
    .b(1'b0),
    .c(al_4090ecdb),
    .o({al_b1c2c144,al_5a529b34[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_21a6a0d7 (
    .a(al_92abc73b[8]),
    .b(1'b1),
    .c(al_b1c2c144),
    .o({al_60d662e6,al_5a529b34[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7610b14 (
    .a(al_92abc73b[9]),
    .b(1'b0),
    .c(al_60d662e6),
    .o({al_687e23a0,al_5a529b34[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d7020d00 (
    .a(al_92abc73b[10]),
    .b(1'b1),
    .c(al_687e23a0),
    .o({al_b5c4be4e,al_5a529b34[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_91d16e11 (
    .a(al_92abc73b[11]),
    .b(1'b0),
    .c(al_b5c4be4e),
    .o({al_f1e4a7a7,al_5a529b34[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b704ba29 (
    .a(al_92abc73b[12]),
    .b(1'b1),
    .c(al_f1e4a7a7),
    .o({al_e2931770,al_5a529b34[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8fcb7c9f (
    .a(al_92abc73b[13]),
    .b(1'b0),
    .c(al_e2931770),
    .o({al_4821ff7f,al_5a529b34[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8ddfc287 (
    .a(al_92abc73b[14]),
    .b(1'b1),
    .c(al_4821ff7f),
    .o({al_712165e6,al_5a529b34[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7402f60d (
    .a(al_92abc73b[15]),
    .b(1'b1),
    .c(al_712165e6),
    .o({al_1749b8de,al_5a529b34[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_417a7a98 (
    .a(al_92abc73b[16]),
    .b(1'b1),
    .c(al_1749b8de),
    .o({al_593536de,al_5a529b34[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_35dea101 (
    .a(al_92abc73b[17]),
    .b(1'b0),
    .c(al_593536de),
    .o({al_8f6c5547,al_5a529b34[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f71f03b6 (
    .a(al_92abc73b[18]),
    .b(1'b1),
    .c(al_8f6c5547),
    .o({al_ff178429,al_5a529b34[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_baac7215 (
    .a(al_92abc73b[19]),
    .b(1'b0),
    .c(al_ff178429),
    .o({al_a46cb2d7,al_5a529b34[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_98dc5fa4 (
    .a(al_92abc73b[20]),
    .b(1'b0),
    .c(al_a46cb2d7),
    .o({al_4e7e9688,al_5a529b34[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e2846a7f (
    .c(al_4e7e9688),
    .o({open_n22,al_5a529b34[20]}));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_fed664a1 (
    .a(al_9ea00fd2),
    .b(num[0]),
    .o(al_6d90eb23[0]));
  AL_MAP_LUT6 #(
    .EQN("(D*~((E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B))*~(A)+D*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*~(A)+~(D)*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*A+D*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*A)"),
    .INIT(64'h7f2a5d0877225500))
    al_98ca4f81 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(al_45db9cb5),
    .d(num[10]),
    .e(num[6]),
    .f(num[2]),
    .o(al_e75a278b));
  AL_MAP_LUT6 #(
    .EQN("(D*~((E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B))*~(A)+D*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*~(A)+~(D)*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*A+D*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*A)"),
    .INIT(64'h7f2a5d0877225500))
    al_61ad8985 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(al_45db9cb5),
    .d(num[11]),
    .e(num[7]),
    .f(num[3]),
    .o(al_57322515));
  AL_MAP_LUT5 #(
    .EQN("(C*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(A)+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)+~(C)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A)"),
    .INIT(32'hfad87250))
    al_6e5744d1 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[12]),
    .d(num[8]),
    .e(num[4]),
    .o(al_e013aab4));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h7430))
    al_980ac878 (
    .a(al_f7b167),
    .b(al_4fb683a3),
    .c(al_e013aab4),
    .d(num[0]),
    .o(al_db63ae90));
  AL_MAP_LUT5 #(
    .EQN("(C*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(A)+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)+~(C)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A)"),
    .INIT(32'hfad87250))
    al_61a44992 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[13]),
    .d(num[9]),
    .e(num[5]),
    .o(al_304d439a));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h7430))
    al_2a78820c (
    .a(al_f7b167),
    .b(al_4fb683a3),
    .c(al_304d439a),
    .d(num[1]),
    .o(al_8bf09624));
  AL_MAP_LUT5 #(
    .EQN("(C*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(A)+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)+~(C)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A)"),
    .INIT(32'hfad87250))
    al_dd57d58d (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[14]),
    .d(num[10]),
    .e(num[6]),
    .o(al_7adb5007));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h7430))
    al_2b7a9f9f (
    .a(al_f7b167),
    .b(al_4fb683a3),
    .c(al_7adb5007),
    .d(num[2]),
    .o(al_6979d612));
  AL_MAP_LUT5 #(
    .EQN("(C*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(A)+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)+~(C)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A)"),
    .INIT(32'hfad87250))
    al_467d28c (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[15]),
    .d(num[11]),
    .e(num[7]),
    .o(al_d5ae2d7f));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h7430))
    al_ab8ccbfc (
    .a(al_f7b167),
    .b(al_4fb683a3),
    .c(al_d5ae2d7f),
    .d(num[3]),
    .o(al_696d4179));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_526de7d8 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(al_36c58aac),
    .d(al_45db9cb5),
    .o(al_f7b167));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_f7f2b4f (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(al_45db9cb5),
    .o(al_4fb683a3));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_3027f931 (
    .a(num[4]),
    .b(num[3]),
    .c(num[2]),
    .d(num[1]),
    .o(al_8c06569d));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_462250c7 (
    .a(al_36c58aac),
    .b(al_8c06569d),
    .o(al_5c9f255f));
  AL_MAP_LUT5 #(
    .EQN("(C*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(A)+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)+~(C)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A+C*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A)"),
    .INIT(32'hfad87250))
    al_46b4dc8c (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[16]),
    .d(num[12]),
    .e(num[8]),
    .o(al_6c0808));
  AL_MAP_LUT6 #(
    .EQN("(D*~((~C*(E*~(F)*~(A)+E*F*~(A)+~(E)*F*A+E*F*A)))*~(B)+D*(~C*(E*~(F)*~(A)+E*F*~(A)+~(E)*F*A+E*F*A))*~(B)+~(D)*(~C*(E*~(F)*~(A)+E*F*~(A)+~(E)*F*A+E*F*A))*B+D*(~C*(E*~(F)*~(A)+E*F*~(A)+~(E)*F*A+E*F*A))*B)"),
    .INIT(64'h3f0c3b0837043300))
    al_86cdbbd (
    .a(al_f7b167),
    .b(al_4fb683a3),
    .c(al_5c9f255f),
    .d(al_6c0808),
    .e(num[4]),
    .f(num[0]),
    .o(al_ae3fe1e5));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_a72e2d94 (
    .a(num[20]),
    .b(num[19]),
    .c(num[18]),
    .d(num[17]),
    .o(al_9ea00fd2));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_f901857b (
    .a(num[16]),
    .b(num[15]),
    .c(num[14]),
    .d(num[13]),
    .o(al_1823807d));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_7038c323 (
    .a(num[8]),
    .b(num[7]),
    .c(num[6]),
    .d(num[5]),
    .o(al_36c58aac));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_3e240b47 (
    .a(num[12]),
    .b(num[11]),
    .c(num[10]),
    .d(num[9]),
    .o(al_45db9cb5));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_cfcdbc2b (
    .a(al_9ea00fd2),
    .b(num[1]),
    .o(al_6d90eb23[1]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_e70474fa (
    .a(al_36c58aac),
    .b(num[8]),
    .c(num[4]),
    .o(al_c3ad1f75));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfaf87270))
    al_da94f4e7 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[20]),
    .d(num[16]),
    .e(num[12]),
    .o(al_788d5b83));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(A*~(C*~(E*B))))"),
    .INIT(32'hff8aff0a))
    al_fada030d (
    .a(al_4fb683a3),
    .b(al_5c9f255f),
    .c(al_c3ad1f75),
    .d(al_788d5b83),
    .e(num[0]),
    .o(al_a980305));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_949fb34f (
    .a(al_9ea00fd2),
    .b(num[2]),
    .o(al_6d90eb23[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_5b5e508b (
    .a(al_9ea00fd2),
    .b(num[3]),
    .o(al_6d90eb23[3]));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    .INIT(16'h7250))
    al_b2c6509f (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[4]),
    .d(num[0]),
    .o(al_6d90eb23[4]));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    .INIT(16'h7250))
    al_6baab633 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[5]),
    .d(num[1]),
    .o(al_6d90eb23[5]));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    .INIT(16'h7250))
    al_1b248346 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[6]),
    .d(num[2]),
    .o(al_6d90eb23[6]));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    .INIT(16'h7250))
    al_d60c418b (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[7]),
    .d(num[3]),
    .o(al_6d90eb23[7]));
  AL_MAP_LUT6 #(
    .EQN("(D*~((E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B))*~(A)+D*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*~(A)+~(D)*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*A+D*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*A)"),
    .INIT(64'h7f2a5d0877225500))
    al_42edd67a (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(al_45db9cb5),
    .d(num[8]),
    .e(num[4]),
    .f(num[0]),
    .o(al_a2611309));
  AL_MAP_LUT6 #(
    .EQN("(D*~((E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B))*~(A)+D*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*~(A)+~(D)*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*A+D*(E*~((F*~C))*~(B)+E*(F*~C)*~(B)+~(E)*(F*~C)*B+E*(F*~C)*B)*A)"),
    .INIT(64'h7f2a5d0877225500))
    al_efc72dd1 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(al_45db9cb5),
    .d(num[9]),
    .e(num[5]),
    .f(num[1]),
    .o(al_3261239f));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(A*~(~D*~(E*B))))"),
    .INIT(32'h0507050f))
    al_eb0bc97b (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[17]),
    .d(num[13]),
    .e(num[9]),
    .o(al_a67b2030));
  AL_MAP_LUT5 #(
    .EQN("(~C*~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*~(B)+~C*(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(B)+~(~C)*(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B+~C*(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*B)"),
    .INIT(32'hcf8b4703))
    al_56d8554b (
    .a(al_f7b167),
    .b(al_4fb683a3),
    .c(al_a67b2030),
    .d(num[5]),
    .e(num[1]),
    .o(al_3123bab1));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(A*~(~D*~(E*B))))"),
    .INIT(32'h0507050f))
    al_90411537 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[18]),
    .d(num[14]),
    .e(num[10]),
    .o(al_8563d1ec));
  AL_MAP_LUT5 #(
    .EQN("~(C*~((D*B)*~(E)*~(A)+(D*B)*E*~(A)+~((D*B))*E*A+(D*B)*E*A))"),
    .INIT(32'hefaf4f0f))
    al_875d7745 (
    .a(al_f7b167),
    .b(al_4fb683a3),
    .c(al_8563d1ec),
    .d(num[6]),
    .e(num[2]),
    .o(al_500d0cf0));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(A*~(~D*~(E*B))))"),
    .INIT(32'h0507050f))
    al_2ef3f387 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(num[19]),
    .d(num[15]),
    .e(num[11]),
    .o(al_fa86226a));
  AL_MAP_LUT5 #(
    .EQN("~(C*~((D*B)*~(E)*~(A)+(D*B)*E*~(A)+~((D*B))*E*A+(D*B)*E*A))"),
    .INIT(32'hefaf4f0f))
    al_5bd2ddb8 (
    .a(al_f7b167),
    .b(al_4fb683a3),
    .c(al_fa86226a),
    .d(num[7]),
    .e(num[3]),
    .o(al_6b3505b5));
  AL_DFF_X al_f54ca955 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6d90eb23[0]),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[0]));
  AL_DFF_X al_2d8af2a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3261239f),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[9]));
  AL_DFF_X al_7a6b8f23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e75a278b),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[10]));
  AL_DFF_X al_66d71082 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57322515),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[11]));
  AL_DFF_X al_90d6e5ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_db63ae90),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[12]));
  AL_DFF_X al_adda3d2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8bf09624),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[13]));
  AL_DFF_X al_4ed8ea65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6979d612),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[14]));
  AL_DFF_X al_40cc5e94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_696d4179),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[15]));
  AL_DFF_X al_6ad454ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ae3fe1e5),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[16]));
  AL_DFF_X al_854e98e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3123bab1),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[17]));
  AL_DFF_X al_2794869c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_500d0cf0),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[18]));
  AL_DFF_X al_fc3f0329 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6d90eb23[1]),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[1]));
  AL_DFF_X al_d88977fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6b3505b5),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[19]));
  AL_DFF_X al_70d1cf85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a980305),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[20]));
  AL_DFF_X al_48d95f6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6d90eb23[2]),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[2]));
  AL_DFF_X al_d4f67b5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6d90eb23[3]),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[3]));
  AL_DFF_X al_231a0942 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6d90eb23[4]),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[4]));
  AL_DFF_X al_65a74cf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6d90eb23[5]),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[5]));
  AL_DFF_X al_6bef8e4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6d90eb23[6]),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[6]));
  AL_DFF_X al_333e0024 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6d90eb23[7]),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[7]));
  AL_DFF_X al_579266e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a2611309),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_92abc73b[8]));
  AL_DFF_X al_35b11324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_de41ded2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(done));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*C*D)"),
    .INIT(16'h1008))
    al_e0d16814 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_fa2e23e1));
  AL_DFF_X al_60e499fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa2e23e1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a7063677));
  AL_DFF_X al_947706c1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_337720e7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b029b709[0]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'ha0b4))
    al_d780acdb (
    .a(al_a7063677),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_803879c7),
    .o(al_82338500));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*(C*B)*~(D)*~(E)+~(A)*~((C*B))*D*~(E)+A*~((C*B))*D*~(E)+A*(C*B)*D*~(E)+A*~((C*B))*D*E+A*(C*B)*D*E)"),
    .INIT(32'haa00bf40))
    al_6533eb33 (
    .a(al_a7063677),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_b029b709[2]),
    .e(al_803879c7),
    .o(al_5669eee7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~((~E*~D*~C))*~(F)+A*B*~((~E*~D*~C))*~(F)+A*B*(~E*~D*~C)*~(F)+~(A)*~(B)*~((~E*~D*~C))*F+~(A)*B*~((~E*~D*~C))*F+A*B*~((~E*~D*~C))*F+~(A)*~(B)*(~E*~D*~C)*F+~(A)*B*(~E*~D*~C)*F+A*B*(~E*~D*~C)*F)"),
    .INIT(64'hdddddddd99999998))
    al_2e877577 (
    .a(al_a7063677),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .f(al_803879c7),
    .o(al_337720e7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*(D*C*B)*~(E)*~(F)+~(A)*~((D*C*B))*E*~(F)+A*~((D*C*B))*E*~(F)+A*(D*C*B)*E*~(F)+A*~((D*C*B))*E*F+A*(D*C*B)*E*F)"),
    .INIT(64'haaaa0000bfff4000))
    al_61a377 (
    .a(al_a7063677),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .f(al_803879c7),
    .o(al_653faf9));
  AL_DFF_X al_5a36a3e9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_82338500),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b029b709[1]));
  AL_DFF_X al_75690eae (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5669eee7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b029b709[2]));
  AL_DFF_X al_67ff022a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_653faf9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b029b709[3]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*~A)"),
    .INIT(32'h00400000))
    al_9830e993 (
    .a(done),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_de41ded2));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_5dd70419 (
    .a(al_de41ded2),
    .b(al_3127e1e8),
    .o(al_c21a53a9[0]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B*~(D*~(~E*C))))"),
    .INIT(32'haa222a22))
    al_e735fd14 (
    .a(al_9ea00fd2),
    .b(al_1823807d),
    .c(al_36c58aac),
    .d(al_45db9cb5),
    .e(al_8c06569d),
    .o(al_338a517[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_574498d2 (
    .a(al_f7b167),
    .b(al_9ea00fd2),
    .c(al_1823807d),
    .o(al_338a517[3]));
  AL_DFF_X al_2adcb2b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_338a517[2]),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e01c36e7[2]));
  AL_DFF_X al_f5c8b177 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_338a517[3]),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e01c36e7[3]));
  AL_DFF_X al_b20c4183 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7b167),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e01c36e7[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_befd69b (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[0]),
    .d(al_16357ce4[2]),
    .e(al_16357ce4[4]),
    .f(al_16357ce4[6]),
    .o(al_54282d1f));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    al_b21f26a0 (
    .a(al_a6672972),
    .b(al_54282d1f),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_b859d315 (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[10]),
    .d(al_16357ce4[12]),
    .e(al_16357ce4[14]),
    .f(al_16357ce4[16]),
    .o(al_3dc3e1bb));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'h003a))
    al_a3b1e637 (
    .a(al_3dc3e1bb),
    .b(al_e1b97ac),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[10]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_42c66aac (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[11]),
    .d(al_16357ce4[13]),
    .e(al_16357ce4[15]),
    .f(al_16357ce4[17]),
    .o(al_fdf9855e));
  AL_MAP_LUT5 #(
    .EQN("(~E*(A*~((~C*B))*~(D)+A*(~C*B)*~(D)+~(A)*(~C*B)*D+A*(~C*B)*D))"),
    .INIT(32'h00000caa))
    al_d0e788cf (
    .a(al_fdf9855e),
    .b(al_f0c918f2),
    .c(al_e01c36e7[3]),
    .d(al_e01c36e7[4]),
    .e(al_3127e1e8),
    .o(al_6de4c23f[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_426b6a39 (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[12]),
    .d(al_16357ce4[14]),
    .e(al_16357ce4[16]),
    .f(al_16357ce4[18]),
    .o(al_83c825e4));
  AL_MAP_LUT5 #(
    .EQN("(~E*(A*~((~C*B))*~(D)+A*(~C*B)*~(D)+~(A)*(~C*B)*D+A*(~C*B)*D))"),
    .INIT(32'h00000caa))
    al_a47e1df2 (
    .a(al_83c825e4),
    .b(al_f3539fe0),
    .c(al_e01c36e7[3]),
    .d(al_e01c36e7[4]),
    .e(al_3127e1e8),
    .o(al_6de4c23f[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_f4ad6f5 (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[13]),
    .d(al_16357ce4[15]),
    .e(al_16357ce4[17]),
    .f(al_16357ce4[19]),
    .o(al_a67e0f03));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~((E*~C*~B))*~(D)+A*(E*~C*~B)*~(D)+~(A)*(E*~C*~B)*D+A*(E*~C*~B)*D))"),
    .INIT(64'h0000000003aa00aa))
    al_12bfc72d (
    .a(al_a67e0f03),
    .b(al_e01c36e7[2]),
    .c(al_e01c36e7[3]),
    .d(al_e01c36e7[4]),
    .e(al_16357ce4[21]),
    .f(al_3127e1e8),
    .o(al_6de4c23f[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_4fd9f712 (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[14]),
    .d(al_16357ce4[16]),
    .e(al_16357ce4[18]),
    .f(al_16357ce4[20]),
    .o(al_a60487f4));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~((E*~C*~B))*~(D)+A*(E*~C*~B)*~(D)+~(A)*(E*~C*~B)*D+A*(E*~C*~B)*D))"),
    .INIT(64'h0000000003aa00aa))
    al_c66921c3 (
    .a(al_a60487f4),
    .b(al_e01c36e7[2]),
    .c(al_e01c36e7[3]),
    .d(al_e01c36e7[4]),
    .e(al_16357ce4[22]),
    .f(al_3127e1e8),
    .o(al_6de4c23f[14]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)*~(C)+(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*~(C)+~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*A*C+(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*C)"),
    .INIT(32'hafaca3a0))
    al_71315719 (
    .a(al_f0c918f2),
    .b(al_e01c36e7[2]),
    .c(al_e01c36e7[3]),
    .d(al_16357ce4[15]),
    .e(al_16357ce4[17]),
    .o(al_dd9cb274));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_36ccc141 (
    .a(al_dd9cb274),
    .b(al_91a73912),
    .o(al_6de4c23f[15]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)*~(C)+(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*~(C)+~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*A*C+(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*C)"),
    .INIT(32'hafaca3a0))
    al_8df200b9 (
    .a(al_f3539fe0),
    .b(al_e01c36e7[2]),
    .c(al_e01c36e7[3]),
    .d(al_16357ce4[16]),
    .e(al_16357ce4[18]),
    .o(al_b050724b));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_3630bbb (
    .a(al_b050724b),
    .b(al_91a73912),
    .o(al_6de4c23f[16]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h89abcdef))
    al_8131fcab (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[17]),
    .d(al_16357ce4[19]),
    .e(al_16357ce4[21]),
    .o(al_8b1fe6d5));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_3c3671b6 (
    .a(al_91a73912),
    .b(al_8b1fe6d5),
    .o(al_6de4c23f[17]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h89abcdef))
    al_5b102fc8 (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[18]),
    .d(al_16357ce4[20]),
    .e(al_16357ce4[22]),
    .o(al_e1b97ac));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_93f4d712 (
    .a(al_91a73912),
    .b(al_e1b97ac),
    .o(al_6de4c23f[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2f99ab87 (
    .a(al_e01c36e7[2]),
    .b(al_16357ce4[19]),
    .c(al_16357ce4[21]),
    .o(al_f0c918f2));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_1ba575ec (
    .a(al_91a73912),
    .b(al_f0c918f2),
    .c(al_e01c36e7[3]),
    .o(al_6de4c23f[19]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_d4daf104 (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[1]),
    .d(al_16357ce4[3]),
    .e(al_16357ce4[5]),
    .f(al_16357ce4[7]),
    .o(al_d3758072));
  AL_MAP_LUT4 #(
    .EQN("(~D*(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h00a3))
    al_4337f44 (
    .a(al_15a841b9),
    .b(al_d3758072),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_891f73c0 (
    .a(al_e01c36e7[4]),
    .b(al_3127e1e8),
    .o(al_91a73912));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_737dfff6 (
    .a(al_e01c36e7[2]),
    .b(al_16357ce4[20]),
    .c(al_16357ce4[22]),
    .o(al_f3539fe0));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_f6e3957 (
    .a(al_91a73912),
    .b(al_f3539fe0),
    .c(al_e01c36e7[3]),
    .o(al_6de4c23f[20]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_636cae6d (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[2]),
    .d(al_16357ce4[4]),
    .e(al_16357ce4[6]),
    .f(al_16357ce4[8]),
    .o(al_75977872));
  AL_MAP_LUT4 #(
    .EQN("(~D*(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h00a3))
    al_184544af (
    .a(al_3dc3e1bb),
    .b(al_75977872),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_c38f30d1 (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[3]),
    .d(al_16357ce4[5]),
    .e(al_16357ce4[7]),
    .f(al_16357ce4[9]),
    .o(al_76d214f0));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    al_19c312a2 (
    .a(al_fdf9855e),
    .b(al_76d214f0),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_67fa2b5d (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[4]),
    .d(al_16357ce4[6]),
    .e(al_16357ce4[8]),
    .f(al_16357ce4[10]),
    .o(al_6067595f));
  AL_MAP_LUT4 #(
    .EQN("(~D*(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h00a3))
    al_b978afeb (
    .a(al_83c825e4),
    .b(al_6067595f),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_1e84725 (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[5]),
    .d(al_16357ce4[7]),
    .e(al_16357ce4[9]),
    .f(al_16357ce4[11]),
    .o(al_babeab3));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    al_2cc7f562 (
    .a(al_a67e0f03),
    .b(al_babeab3),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_17dd233f (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[6]),
    .d(al_16357ce4[8]),
    .e(al_16357ce4[10]),
    .f(al_16357ce4[12]),
    .o(al_ab2fd291));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    al_67ea44e8 (
    .a(al_a60487f4),
    .b(al_ab2fd291),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_baa3bf0f (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[7]),
    .d(al_16357ce4[9]),
    .e(al_16357ce4[11]),
    .f(al_16357ce4[13]),
    .o(al_2b66b96f));
  AL_MAP_LUT4 #(
    .EQN("(~D*(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h00a3))
    al_93388a29 (
    .a(al_dd9cb274),
    .b(al_2b66b96f),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_c262e922 (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[8]),
    .d(al_16357ce4[10]),
    .e(al_16357ce4[12]),
    .f(al_16357ce4[14]),
    .o(al_a6672972));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    al_ea54a76 (
    .a(al_b050724b),
    .b(al_a6672972),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_b2eaa791 (
    .a(al_e01c36e7[2]),
    .b(al_e01c36e7[3]),
    .c(al_16357ce4[9]),
    .d(al_16357ce4[11]),
    .e(al_16357ce4[13]),
    .f(al_16357ce4[15]),
    .o(al_15a841b9));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'h003a))
    al_15a467f6 (
    .a(al_15a841b9),
    .b(al_8b1fe6d5),
    .c(al_e01c36e7[4]),
    .d(al_3127e1e8),
    .o(al_6de4c23f[9]));
  AL_DFF_X al_1e3b351c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[0]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[0]));
  AL_DFF_X al_5c59aaac (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[9]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[9]));
  AL_DFF_X al_3e347a3e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[10]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[10]));
  AL_DFF_X al_c5fe0851 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[11]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[11]));
  AL_DFF_X al_c8ed733f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[12]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[12]));
  AL_DFF_X al_b53f7182 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[13]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[13]));
  AL_DFF_X al_673b2e41 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[14]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[14]));
  AL_DFF_X al_5fba0afb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[15]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[15]));
  AL_DFF_X al_2bceeb5b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[16]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[16]));
  AL_DFF_X al_7a8e17c3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[17]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[17]));
  AL_DFF_X al_46a26753 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[18]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[18]));
  AL_DFF_X al_9674742 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[1]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[1]));
  AL_DFF_X al_98940337 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[19]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[19]));
  AL_DFF_X al_56210d16 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[20]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[20]));
  AL_DFF_X al_5adc81b0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[2]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[2]));
  AL_DFF_X al_992288cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[3]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[3]));
  AL_DFF_X al_bd7304a0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[4]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[4]));
  AL_DFF_X al_d7824021 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[5]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[5]));
  AL_DFF_X al_8174d8f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[6]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[6]));
  AL_DFF_X al_18798991 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[7]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[7]));
  AL_DFF_X al_22e0cf5c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6de4c23f[8]),
    .en(al_c21a53a9[0]),
    .sr(1'b0),
    .ss(1'b0),
    .q(sqrt[8]));
  AL_DFF_X al_dce734fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(start),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_803879c7));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b9c8457 (
    .a(al_16357ce4[7]),
    .b(al_19b5d2a2[7]),
    .c(al_dc44be48),
    .o({al_d8dd00e3,al_8ff04cfd[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e613dd7 (
    .a(al_16357ce4[8]),
    .b(al_19b5d2a2[8]),
    .c(al_d8dd00e3),
    .o({al_a0bad8f5,al_8ff04cfd[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27c8842d (
    .a(al_16357ce4[9]),
    .b(al_19b5d2a2[9]),
    .c(al_a0bad8f5),
    .o({al_c93e73fa,al_8ff04cfd[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_462a01f1 (
    .a(al_16357ce4[10]),
    .b(al_19b5d2a2[10]),
    .c(al_c93e73fa),
    .o({al_6ea85cef,al_8ff04cfd[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b3bce39 (
    .a(al_16357ce4[11]),
    .b(al_19b5d2a2[11]),
    .c(al_6ea85cef),
    .o({al_52616de9,al_8ff04cfd[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f829bb24 (
    .a(al_16357ce4[12]),
    .b(al_19b5d2a2[12]),
    .c(al_52616de9),
    .o({al_ec1119c9,al_8ff04cfd[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc29264d (
    .a(al_16357ce4[13]),
    .b(al_19b5d2a2[13]),
    .c(al_ec1119c9),
    .o({al_77f3553d,al_8ff04cfd[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee4a1d93 (
    .a(al_16357ce4[14]),
    .b(al_19b5d2a2[14]),
    .c(al_77f3553d),
    .o({al_6299424f,al_8ff04cfd[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_154312aa (
    .a(al_16357ce4[15]),
    .b(al_19b5d2a2[15]),
    .c(al_6299424f),
    .o({al_ea5880d3,al_8ff04cfd[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17566e78 (
    .a(al_16357ce4[16]),
    .b(al_19b5d2a2[16]),
    .c(al_ea5880d3),
    .o({al_bbe9aae2,al_8ff04cfd[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f5224f5b (
    .a(1'b0),
    .o({al_ae0a6293,open_n25}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_38657e34 (
    .a(al_16357ce4[17]),
    .b(al_19b5d2a2[17]),
    .c(al_bbe9aae2),
    .o({al_d9ef6091,al_8ff04cfd[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bbcbdbe (
    .a(al_16357ce4[18]),
    .b(al_19b5d2a2[18]),
    .c(al_d9ef6091),
    .o({al_7109a3cd,al_8ff04cfd[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_216ec453 (
    .a(al_16357ce4[19]),
    .b(al_19b5d2a2[19]),
    .c(al_7109a3cd),
    .o({al_f1bac0a6,al_8ff04cfd[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c943a4d2 (
    .a(al_16357ce4[20]),
    .b(al_19b5d2a2[20]),
    .c(al_f1bac0a6),
    .o({al_61c118b2,al_8ff04cfd[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_920ee641 (
    .a(al_16357ce4[21]),
    .b(al_19b5d2a2[21]),
    .c(al_61c118b2),
    .o({al_9bb03b7,al_8ff04cfd[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e359bb16 (
    .a(al_16357ce4[22]),
    .b(al_19b5d2a2[21]),
    .c(al_9bb03b7),
    .o({open_n26,al_8ff04cfd[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e6e3dfcf (
    .a(al_16357ce4[0]),
    .b(al_19b5d2a2[0]),
    .c(al_ae0a6293),
    .o({al_d07a623a,al_8ff04cfd[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68abff86 (
    .a(al_16357ce4[1]),
    .b(al_19b5d2a2[1]),
    .c(al_d07a623a),
    .o({al_126bbf82,al_8ff04cfd[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8de058bd (
    .a(al_16357ce4[2]),
    .b(al_19b5d2a2[2]),
    .c(al_126bbf82),
    .o({al_1aac3445,al_8ff04cfd[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbd4c846 (
    .a(al_16357ce4[3]),
    .b(al_19b5d2a2[3]),
    .c(al_1aac3445),
    .o({al_f5516224,al_8ff04cfd[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_222b6767 (
    .a(al_16357ce4[4]),
    .b(al_19b5d2a2[4]),
    .c(al_f5516224),
    .o({al_91108e0e,al_8ff04cfd[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c7fbfa5 (
    .a(al_16357ce4[5]),
    .b(al_19b5d2a2[5]),
    .c(al_91108e0e),
    .o({al_a4e1781b,al_8ff04cfd[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd218d47 (
    .a(al_16357ce4[6]),
    .b(al_19b5d2a2[6]),
    .c(al_a4e1781b),
    .o({al_dc44be48,al_8ff04cfd[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4dfdc771 (
    .a(al_da03ca6b[7]),
    .b(al_7b2fe207[7]),
    .c(al_5d663e44),
    .o({al_27011e73,al_de90ce1b[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e93dcd8b (
    .a(al_da03ca6b[8]),
    .b(al_7b2fe207[8]),
    .c(al_27011e73),
    .o({al_4c0f5956,al_de90ce1b[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2f94769 (
    .a(al_da03ca6b[9]),
    .b(al_7b2fe207[9]),
    .c(al_4c0f5956),
    .o({al_e0589574,al_de90ce1b[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_18f640ef (
    .a(al_da03ca6b[10]),
    .b(al_7b2fe207[10]),
    .c(al_e0589574),
    .o({al_12f8fb3c,al_de90ce1b[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86ec8670 (
    .a(al_da03ca6b[11]),
    .b(al_7b2fe207[11]),
    .c(al_12f8fb3c),
    .o({al_3c4a6475,al_de90ce1b[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6df03772 (
    .a(al_da03ca6b[12]),
    .b(al_7b2fe207[12]),
    .c(al_3c4a6475),
    .o({al_9fa575eb,al_de90ce1b[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_45f02cda (
    .a(al_da03ca6b[13]),
    .b(al_7b2fe207[13]),
    .c(al_9fa575eb),
    .o({al_d3327d96,al_de90ce1b[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f6b2c7c5 (
    .a(al_da03ca6b[14]),
    .b(al_7b2fe207[14]),
    .c(al_d3327d96),
    .o({al_412f61d0,al_de90ce1b[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86f06d29 (
    .a(al_da03ca6b[15]),
    .b(al_7b2fe207[15]),
    .c(al_412f61d0),
    .o({al_3b62f46f,al_de90ce1b[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff64c9f9 (
    .a(al_da03ca6b[16]),
    .b(al_7b2fe207[16]),
    .c(al_3b62f46f),
    .o({al_5d141531,al_de90ce1b[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_6219435f (
    .a(1'b0),
    .o({al_d6d4ff9e,open_n29}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_689e06a4 (
    .a(al_da03ca6b[17]),
    .b(al_7b2fe207[17]),
    .c(al_5d141531),
    .o({al_67aa9deb,al_de90ce1b[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a011db00 (
    .a(al_da03ca6b[18]),
    .b(al_7b2fe207[18]),
    .c(al_67aa9deb),
    .o({al_3697e743,al_de90ce1b[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ebcca0b3 (
    .a(al_da03ca6b[19]),
    .b(al_7b2fe207[19]),
    .c(al_3697e743),
    .o({al_3d62c9fe,al_de90ce1b[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b00f8a2c (
    .a(al_da03ca6b[20]),
    .b(al_7b2fe207[20]),
    .c(al_3d62c9fe),
    .o({al_81a11f5a,al_de90ce1b[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_67573096 (
    .a(al_da03ca6b[21]),
    .b(al_7b2fe207[21]),
    .c(al_81a11f5a),
    .o({al_461d7931,al_de90ce1b[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a4bf0f3d (
    .a(al_da03ca6b[22]),
    .b(al_7b2fe207[21]),
    .c(al_461d7931),
    .o({open_n30,al_de90ce1b[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9173b3c2 (
    .a(al_da03ca6b[0]),
    .b(al_7b2fe207[0]),
    .c(al_d6d4ff9e),
    .o({al_b6ba68ca,al_de90ce1b[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1e14f1c1 (
    .a(al_da03ca6b[1]),
    .b(al_7b2fe207[1]),
    .c(al_b6ba68ca),
    .o({al_3c3af6b1,al_de90ce1b[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b174dbc (
    .a(al_da03ca6b[2]),
    .b(al_7b2fe207[2]),
    .c(al_3c3af6b1),
    .o({al_c7e7c580,al_de90ce1b[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6657a45b (
    .a(al_da03ca6b[3]),
    .b(al_7b2fe207[3]),
    .c(al_c7e7c580),
    .o({al_a93520ae,al_de90ce1b[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17e08140 (
    .a(al_da03ca6b[4]),
    .b(al_7b2fe207[4]),
    .c(al_a93520ae),
    .o({al_81c04c9c,al_de90ce1b[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e94e10ff (
    .a(al_da03ca6b[5]),
    .b(al_7b2fe207[5]),
    .c(al_81c04c9c),
    .o({al_f584a17a,al_de90ce1b[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_440a3abe (
    .a(al_da03ca6b[6]),
    .b(al_7b2fe207[6]),
    .c(al_f584a17a),
    .o({al_5d663e44,al_de90ce1b[6]}));
  AL_MAP_LUT5 #(
    .EQN("((D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*~(B)*~(C)+(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*B*~(C)+~((D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E))*B*C+(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*B*C)"),
    .INIT(32'hcacacfc0))
    al_362811ad (
    .a(al_d65643ad[0]),
    .b(al_92abc73b[0]),
    .c(al_803879c7),
    .d(al_8ff04cfd[0]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[0]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_ac6014fb (
    .a(al_378a1ee4[9]),
    .b(al_d65643ad[10]),
    .c(al_803879c7),
    .d(al_8ff04cfd[10]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[10]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_64f81a80 (
    .a(al_378a1ee4[10]),
    .b(al_d65643ad[11]),
    .c(al_803879c7),
    .d(al_8ff04cfd[11]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[11]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_b89c7a41 (
    .a(al_378a1ee4[11]),
    .b(al_d65643ad[12]),
    .c(al_803879c7),
    .d(al_8ff04cfd[12]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[12]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_2f3cde41 (
    .a(al_378a1ee4[12]),
    .b(al_d65643ad[13]),
    .c(al_803879c7),
    .d(al_8ff04cfd[13]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[13]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_551fb630 (
    .a(al_378a1ee4[13]),
    .b(al_d65643ad[14]),
    .c(al_803879c7),
    .d(al_8ff04cfd[14]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[14]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_5e3f3097 (
    .a(al_378a1ee4[14]),
    .b(al_d65643ad[15]),
    .c(al_803879c7),
    .d(al_8ff04cfd[15]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[15]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_32aabe1b (
    .a(al_378a1ee4[15]),
    .b(al_d65643ad[16]),
    .c(al_803879c7),
    .d(al_8ff04cfd[16]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[16]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_a04b95e6 (
    .a(al_378a1ee4[16]),
    .b(al_d65643ad[17]),
    .c(al_803879c7),
    .d(al_8ff04cfd[17]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[17]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_87c5cb1 (
    .a(al_378a1ee4[17]),
    .b(al_d65643ad[18]),
    .c(al_803879c7),
    .d(al_8ff04cfd[18]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[18]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_c7a1d390 (
    .a(al_378a1ee4[18]),
    .b(al_d65643ad[19]),
    .c(al_803879c7),
    .d(al_8ff04cfd[19]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[19]));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*~(B)*~(C)+~(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*B*~(C)+~(~(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E))*B*C+~(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*B*C)"),
    .INIT(32'h3a3a3f30))
    al_3895a34b (
    .a(al_d65643ad[1]),
    .b(al_92abc73b[1]),
    .c(al_803879c7),
    .d(al_8ff04cfd[1]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[1]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_c2f0948c (
    .a(al_378a1ee4[19]),
    .b(al_d65643ad[20]),
    .c(al_803879c7),
    .d(al_8ff04cfd[20]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[20]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_a2c69e49 (
    .a(al_6f8464f),
    .b(al_d65643ad[21]),
    .c(al_803879c7),
    .d(al_8ff04cfd[21]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[21]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_7045eaf3 (
    .a(al_378a1ee4[1]),
    .b(al_d65643ad[2]),
    .c(al_803879c7),
    .d(al_8ff04cfd[2]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[2]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_74e048af (
    .a(al_378a1ee4[2]),
    .b(al_d65643ad[3]),
    .c(al_803879c7),
    .d(al_8ff04cfd[3]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[3]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_ef2081cf (
    .a(al_378a1ee4[3]),
    .b(al_d65643ad[4]),
    .c(al_803879c7),
    .d(al_8ff04cfd[4]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[4]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_65c4b02d (
    .a(al_378a1ee4[4]),
    .b(al_d65643ad[5]),
    .c(al_803879c7),
    .d(al_8ff04cfd[5]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[5]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_ae0353f1 (
    .a(al_378a1ee4[5]),
    .b(al_d65643ad[6]),
    .c(al_803879c7),
    .d(al_8ff04cfd[6]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[6]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_d2584d4b (
    .a(al_378a1ee4[6]),
    .b(al_d65643ad[7]),
    .c(al_803879c7),
    .d(al_8ff04cfd[7]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[7]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_dea0726d (
    .a(al_378a1ee4[7]),
    .b(al_d65643ad[8]),
    .c(al_803879c7),
    .d(al_8ff04cfd[8]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[8]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'hacacafa0))
    al_fb27239 (
    .a(al_378a1ee4[8]),
    .b(al_d65643ad[9]),
    .c(al_803879c7),
    .d(al_8ff04cfd[9]),
    .e(al_da03ca6b[22]),
    .o(al_f8bbbf13[9]));
  AL_DFF_X al_5cc6d5b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[0]));
  AL_DFF_X al_4db9b8f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[9]));
  AL_DFF_X al_c37f14c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[10]));
  AL_DFF_X al_6d92ed15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[11]));
  AL_DFF_X al_33dde6ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[12]));
  AL_DFF_X al_705369da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[13]));
  AL_DFF_X al_6bccd639 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[14]));
  AL_DFF_X al_2c49574e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[15]));
  AL_DFF_X al_55f26226 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[16]));
  AL_DFF_X al_25dfb10f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[17]));
  AL_DFF_X al_dd7cf631 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[18]));
  AL_DFF_X al_81d45cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[1]));
  AL_DFF_X al_5dda0a3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[19]));
  AL_DFF_X al_e52ef9ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[20]));
  AL_DFF_X al_7131e5c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[21]));
  AL_DFF_X al_1c19e6ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_42fa3115),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[22]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .INIT(16'h2230))
    al_a9c9d151 (
    .a(al_d65643ad[22]),
    .b(al_803879c7),
    .c(al_8ff04cfd[22]),
    .d(al_da03ca6b[22]),
    .o(al_42fa3115));
  AL_DFF_X al_f2c72a20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[2]));
  AL_DFF_X al_348fb3fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[3]));
  AL_DFF_X al_77fefb61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[4]));
  AL_DFF_X al_2e432f53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[5]));
  AL_DFF_X al_b08c3897 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[6]));
  AL_DFF_X al_c9436840 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[7]));
  AL_DFF_X al_9e2095be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8bbbf13[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16357ce4[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_15f604ea (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[0]),
    .d(al_16357ce4[1]),
    .e(al_16357ce4[2]),
    .f(al_16357ce4[3]),
    .o(al_534eeb32));
  AL_MAP_LUT5 #(
    .EQN("((~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)*~(A)*~(E)+(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)*A*~(E)+~((~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D))*A*E+(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)*A*E)"),
    .INIT(32'haaaaf033))
    al_98f28111 (
    .a(al_ded0a164),
    .b(al_534eeb32),
    .c(al_7406b7f),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_7b2fe207[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff0ccaa00f0ccaa))
    al_76ab35c6 (
    .a(al_a65c875a),
    .b(al_da2dd23a),
    .c(al_b2a2e5ce),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .f(al_16357ce4[22]),
    .o(al_7b2fe207[10]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff0ccaa00f0ccaa))
    al_a4b24f0a (
    .a(al_43cf9c51),
    .b(al_312b9047),
    .c(al_fe92b9c9),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .f(al_16357ce4[22]),
    .o(al_7b2fe207[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f6aaef9b (
    .a(al_f3ac4ff4),
    .b(al_462198a),
    .c(al_b029b709[2]),
    .o(al_6bd399c8));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_a23c8cd4 (
    .a(al_1f8ac62a),
    .b(al_b029b709[2]),
    .c(al_16357ce4[22]),
    .o(al_14573418));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_12a219f9 (
    .a(al_6bd399c8),
    .b(al_14573418),
    .c(al_b029b709[3]),
    .o(al_7b2fe207[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_36300d15 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[13]),
    .d(al_16357ce4[14]),
    .e(al_16357ce4[15]),
    .f(al_16357ce4[16]),
    .o(al_fb75ed64));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_304017e7 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[17]),
    .d(al_16357ce4[18]),
    .e(al_16357ce4[19]),
    .f(al_16357ce4[20]),
    .o(al_c9156751));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f172a0e3 (
    .a(al_fb75ed64),
    .b(al_c9156751),
    .c(al_b029b709[2]),
    .o(al_2ec9e601));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((~C*~B*~A))+E*D*~((~C*~B*~A))+~(E)*D*(~C*~B*~A)+E*D*(~C*~B*~A))"),
    .INIT(32'hfffe0100))
    al_ba8904ca (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_b029b709[2]),
    .d(al_16357ce4[21]),
    .e(al_16357ce4[22]),
    .o(al_db11fb22));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e6b06aae (
    .a(al_2ec9e601),
    .b(al_db11fb22),
    .c(al_b029b709[3]),
    .o(al_7b2fe207[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_57cbccd8 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[14]),
    .d(al_16357ce4[15]),
    .e(al_16357ce4[16]),
    .f(al_16357ce4[17]),
    .o(al_da2dd23a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_6392c188 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[18]),
    .d(al_16357ce4[19]),
    .e(al_16357ce4[20]),
    .f(al_16357ce4[21]),
    .o(al_b2a2e5ce));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(E)*~(D)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*~(D)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*E*D+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*D)"),
    .INIT(32'hffca00ca))
    al_a3f1e55f (
    .a(al_da2dd23a),
    .b(al_b2a2e5ce),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .e(al_16357ce4[22]),
    .o(al_7b2fe207[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_c0f098a (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[15]),
    .d(al_16357ce4[16]),
    .e(al_16357ce4[17]),
    .f(al_16357ce4[18]),
    .o(al_312b9047));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_cfa70f8b (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[19]),
    .d(al_16357ce4[20]),
    .e(al_16357ce4[21]),
    .f(al_16357ce4[22]),
    .o(al_fe92b9c9));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(E)*~(D)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*~(D)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*E*D+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*D)"),
    .INIT(32'hffca00ca))
    al_b5132400 (
    .a(al_312b9047),
    .b(al_fe92b9c9),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .e(al_16357ce4[22]),
    .o(al_7b2fe207[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_6a540ef8 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[16]),
    .d(al_16357ce4[17]),
    .e(al_16357ce4[18]),
    .f(al_16357ce4[19]),
    .o(al_462198a));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    al_ff8e5f2c (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[20]),
    .d(al_16357ce4[21]),
    .e(al_16357ce4[22]),
    .o(al_1f8ac62a));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(E)*~(D)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*~(D)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*E*D+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*D)"),
    .INIT(32'hffca00ca))
    al_c39e36de (
    .a(al_462198a),
    .b(al_1f8ac62a),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .e(al_16357ce4[22]),
    .o(al_7b2fe207[16]));
  AL_MAP_LUT6 #(
    .EQN("(A*~((F*~(E)*~((~C*~B))+F*E*~((~C*~B))+~(F)*E*(~C*~B)+F*E*(~C*~B)))*~(D)+A*(F*~(E)*~((~C*~B))+F*E*~((~C*~B))+~(F)*E*(~C*~B)+F*E*(~C*~B))*~(D)+~(A)*(F*~(E)*~((~C*~B))+F*E*~((~C*~B))+~(F)*E*(~C*~B)+F*E*(~C*~B))*D+A*(F*~(E)*~((~C*~B))+F*E*~((~C*~B))+~(F)*E*(~C*~B)+F*E*(~C*~B))*D)"),
    .INIT(64'hffaafcaa03aa00aa))
    al_31ed852e (
    .a(al_c9156751),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_b029b709[2]),
    .e(al_16357ce4[21]),
    .f(al_16357ce4[22]),
    .o(al_c6dd6de));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_6fe5df2d (
    .a(al_c6dd6de),
    .b(al_b029b709[3]),
    .c(al_16357ce4[22]),
    .o(al_7b2fe207[17]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A)*~((~C*~B))+D*A*~((~C*~B))+~(D)*A*(~C*~B)+D*A*(~C*~B))"),
    .INIT(16'hfe02))
    al_517ab28d (
    .a(al_b2a2e5ce),
    .b(al_b029b709[2]),
    .c(al_b029b709[3]),
    .d(al_16357ce4[22]),
    .o(al_7b2fe207[18]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A)*~((~C*~B))+D*A*~((~C*~B))+~(D)*A*(~C*~B)+D*A*(~C*~B))"),
    .INIT(16'hfe02))
    al_e6ca4010 (
    .a(al_fe92b9c9),
    .b(al_b029b709[2]),
    .c(al_b029b709[3]),
    .d(al_16357ce4[22]),
    .o(al_7b2fe207[19]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_8fa46caf (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[1]),
    .d(al_16357ce4[2]),
    .e(al_16357ce4[3]),
    .f(al_16357ce4[4]),
    .o(al_1ea08bcc));
  AL_MAP_LUT5 #(
    .EQN("((~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)*~(A)*~(E)+(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)*A*~(E)+~((~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D))*A*E+(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)*A*E)"),
    .INIT(32'haaaaf033))
    al_41e20a70 (
    .a(al_1e89e993),
    .b(al_1ea08bcc),
    .c(al_b81bed99),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_7b2fe207[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_57eaf2e2 (
    .a(al_14573418),
    .b(al_b029b709[3]),
    .c(al_16357ce4[22]),
    .o(al_7b2fe207[20]));
  AL_MAP_LUT6 #(
    .EQN("(F*~(E)*~((~D*~C*~B*~A))+F*E*~((~D*~C*~B*~A))+~(F)*E*(~D*~C*~B*~A)+F*E*(~D*~C*~B*~A))"),
    .INIT(64'hfffffffe00010000))
    al_81d16c70 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .e(al_16357ce4[21]),
    .f(al_16357ce4[22]),
    .o(al_7b2fe207[21]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_3fea6048 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[2]),
    .d(al_16357ce4[3]),
    .e(al_16357ce4[4]),
    .f(al_16357ce4[5]),
    .o(al_81b0c7fb));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccaaaaff00f0f0))
    al_e542b7a2 (
    .a(al_a65c875a),
    .b(al_da2dd23a),
    .c(al_81b0c7fb),
    .d(al_f33a944d),
    .e(al_b029b709[2]),
    .f(al_b029b709[3]),
    .o(al_7b2fe207[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_9dc84cc8 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[3]),
    .d(al_16357ce4[4]),
    .e(al_16357ce4[5]),
    .f(al_16357ce4[6]),
    .o(al_3896e32f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccaaaaff000f0f))
    al_dbe9321b (
    .a(al_43cf9c51),
    .b(al_312b9047),
    .c(al_3896e32f),
    .d(al_86dcc04b),
    .e(al_b029b709[2]),
    .f(al_b029b709[3]),
    .o(al_7b2fe207[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_4ea0dd64 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[4]),
    .d(al_16357ce4[5]),
    .e(al_16357ce4[6]),
    .f(al_16357ce4[7]),
    .o(al_7406b7f));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(E)+(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(E)+~((C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*E+(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*E)"),
    .INIT(32'haaaaccf0))
    al_488a8738 (
    .a(al_6bd399c8),
    .b(al_68be76e6),
    .c(al_7406b7f),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_7b2fe207[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_66b991b5 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[5]),
    .d(al_16357ce4[6]),
    .e(al_16357ce4[7]),
    .f(al_16357ce4[8]),
    .o(al_b81bed99));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(E)+(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(E)+~((C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*E+(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*E)"),
    .INIT(32'haaaaccf0))
    al_bff6f4c0 (
    .a(al_2ec9e601),
    .b(al_64d5f40e),
    .c(al_b81bed99),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_7b2fe207[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_e8f096bf (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[10]),
    .d(al_16357ce4[11]),
    .e(al_16357ce4[12]),
    .f(al_16357ce4[13]),
    .o(al_a65c875a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_640364b2 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[6]),
    .d(al_16357ce4[7]),
    .e(al_16357ce4[8]),
    .f(al_16357ce4[9]),
    .o(al_f33a944d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00ccccaaaaf0f0))
    al_281296a8 (
    .a(al_a65c875a),
    .b(al_da2dd23a),
    .c(al_f33a944d),
    .d(al_b2a2e5ce),
    .e(al_b029b709[2]),
    .f(al_b029b709[3]),
    .o(al_7b2fe207[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_fc0f7b67 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[11]),
    .d(al_16357ce4[12]),
    .e(al_16357ce4[13]),
    .f(al_16357ce4[14]),
    .o(al_43cf9c51));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_5abcf85 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[7]),
    .d(al_16357ce4[8]),
    .e(al_16357ce4[9]),
    .f(al_16357ce4[10]),
    .o(al_86dcc04b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00ccccaaaaf0f0))
    al_3ae57c40 (
    .a(al_43cf9c51),
    .b(al_312b9047),
    .c(al_86dcc04b),
    .d(al_fe92b9c9),
    .e(al_b029b709[2]),
    .f(al_b029b709[3]),
    .o(al_7b2fe207[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_106815f2 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[8]),
    .d(al_16357ce4[9]),
    .e(al_16357ce4[10]),
    .f(al_16357ce4[11]),
    .o(al_68be76e6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_2a8b36dc (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[12]),
    .d(al_16357ce4[13]),
    .e(al_16357ce4[14]),
    .f(al_16357ce4[15]),
    .o(al_f3ac4ff4));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a889d983 (
    .a(al_68be76e6),
    .b(al_f3ac4ff4),
    .c(al_b029b709[2]),
    .o(al_ded0a164));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E)"),
    .INIT(32'hf0ccaaaa))
    al_a2a62334 (
    .a(al_ded0a164),
    .b(al_462198a),
    .c(al_1f8ac62a),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_7b2fe207[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_3119494e (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_16357ce4[9]),
    .d(al_16357ce4[10]),
    .e(al_16357ce4[11]),
    .f(al_16357ce4[12]),
    .o(al_64d5f40e));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_81a064c6 (
    .a(al_64d5f40e),
    .b(al_fb75ed64),
    .c(al_b029b709[2]),
    .o(al_1e89e993));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_538ce014 (
    .a(al_1e89e993),
    .b(al_c6dd6de),
    .c(al_b029b709[3]),
    .o(al_7b2fe207[9]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*~(B)*~(C)+(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*B*~(C)+~((D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E))*B*C+(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*B*C)"),
    .INIT(32'hcacacfc0))
    al_cdd2d16e (
    .a(al_c968c273[0]),
    .b(al_92abc73b[0]),
    .c(al_803879c7),
    .d(al_de90ce1b[0]),
    .e(al_da03ca6b[22]),
    .o(al_cbee0ff9[0]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_cadb5222 (
    .a(al_c968c273[10]),
    .b(al_803879c7),
    .c(al_de90ce1b[10]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[9]),
    .o(al_cbee0ff9[10]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_ddb9e65f (
    .a(al_c968c273[11]),
    .b(al_803879c7),
    .c(al_de90ce1b[11]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[10]),
    .o(al_cbee0ff9[11]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_179f3a29 (
    .a(al_c968c273[12]),
    .b(al_803879c7),
    .c(al_de90ce1b[12]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[11]),
    .o(al_cbee0ff9[12]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_d34153cd (
    .a(al_c968c273[13]),
    .b(al_803879c7),
    .c(al_de90ce1b[13]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[12]),
    .o(al_cbee0ff9[13]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_9d56ed5f (
    .a(al_c968c273[14]),
    .b(al_803879c7),
    .c(al_de90ce1b[14]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[13]),
    .o(al_cbee0ff9[14]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_5599c2a0 (
    .a(al_c968c273[15]),
    .b(al_803879c7),
    .c(al_de90ce1b[15]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[14]),
    .o(al_cbee0ff9[15]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_c349ca41 (
    .a(al_c968c273[16]),
    .b(al_803879c7),
    .c(al_de90ce1b[16]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[15]),
    .o(al_cbee0ff9[16]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_67e777b3 (
    .a(al_c968c273[17]),
    .b(al_803879c7),
    .c(al_de90ce1b[17]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[16]),
    .o(al_cbee0ff9[17]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_e15b33be (
    .a(al_c968c273[18]),
    .b(al_803879c7),
    .c(al_de90ce1b[18]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[17]),
    .o(al_cbee0ff9[18]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_97159ad6 (
    .a(al_c968c273[19]),
    .b(al_803879c7),
    .c(al_de90ce1b[19]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[18]),
    .o(al_cbee0ff9[19]));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*~(B)*~(C)+~(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*B*~(C)+~(~(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E))*B*C+~(D*~(A)*~(E)+D*A*~(E)+~(D)*A*E+D*A*E)*B*C)"),
    .INIT(32'h3a3a3f30))
    al_46c4d16c (
    .a(al_c968c273[1]),
    .b(al_92abc73b[1]),
    .c(al_803879c7),
    .d(al_de90ce1b[1]),
    .e(al_da03ca6b[22]),
    .o(al_cbee0ff9[1]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_3ed4276 (
    .a(al_c968c273[20]),
    .b(al_803879c7),
    .c(al_de90ce1b[20]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[19]),
    .o(al_cbee0ff9[20]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_d32decf4 (
    .a(al_c968c273[21]),
    .b(al_803879c7),
    .c(al_de90ce1b[21]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[20]),
    .o(al_cbee0ff9[21]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_672c0b83 (
    .a(al_c968c273[22]),
    .b(al_803879c7),
    .c(al_de90ce1b[22]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[20]),
    .o(al_cbee0ff9[22]));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(A)*~(C)+~(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*~(C)+~(~(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*A*C+~(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*A*C)"),
    .INIT(32'h5c5c5f50))
    al_83d653b5 (
    .a(al_378a1ee4[1]),
    .b(al_c968c273[2]),
    .c(al_803879c7),
    .d(al_de90ce1b[2]),
    .e(al_da03ca6b[22]),
    .o(al_cbee0ff9[2]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_f54908c8 (
    .a(al_c968c273[3]),
    .b(al_803879c7),
    .c(al_de90ce1b[3]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[2]),
    .o(al_cbee0ff9[3]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_424fd23 (
    .a(al_c968c273[4]),
    .b(al_803879c7),
    .c(al_de90ce1b[4]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[3]),
    .o(al_cbee0ff9[4]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_19dd6680 (
    .a(al_c968c273[5]),
    .b(al_803879c7),
    .c(al_de90ce1b[5]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[4]),
    .o(al_cbee0ff9[5]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_7b2de1ed (
    .a(al_c968c273[6]),
    .b(al_803879c7),
    .c(al_de90ce1b[6]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[5]),
    .o(al_cbee0ff9[6]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_dcb0ecd0 (
    .a(al_c968c273[7]),
    .b(al_803879c7),
    .c(al_de90ce1b[7]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[6]),
    .o(al_cbee0ff9[7]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_92cffc75 (
    .a(al_c968c273[8]),
    .b(al_803879c7),
    .c(al_de90ce1b[8]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[7]),
    .o(al_cbee0ff9[8]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'heefc2230))
    al_8c388bb4 (
    .a(al_c968c273[9]),
    .b(al_803879c7),
    .c(al_de90ce1b[9]),
    .d(al_da03ca6b[22]),
    .e(al_5a529b34[8]),
    .o(al_cbee0ff9[9]));
  AL_DFF_X al_74ba8a60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[0]));
  AL_DFF_X al_f49fce43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[9]));
  AL_DFF_X al_4d88b3ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[10]));
  AL_DFF_X al_d13bc574 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[11]));
  AL_DFF_X al_a89fe0ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[12]));
  AL_DFF_X al_9ed2d193 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[13]));
  AL_DFF_X al_f5437d35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[14]));
  AL_DFF_X al_c6c91e44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[15]));
  AL_DFF_X al_76397f91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[16]));
  AL_DFF_X al_2b6eb27c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[17]));
  AL_DFF_X al_671aacee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[18]));
  AL_DFF_X al_48ba44c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[1]));
  AL_DFF_X al_19664964 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[19]));
  AL_DFF_X al_76de5bd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[20]));
  AL_DFF_X al_ba1f4c46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[21]));
  AL_DFF_X al_51040d30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[22]));
  AL_DFF_X al_8efe335a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[2]));
  AL_DFF_X al_99e618c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[3]));
  AL_DFF_X al_2b9a84c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[4]));
  AL_DFF_X al_9d25a4d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[5]));
  AL_DFF_X al_5564df4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[6]));
  AL_DFF_X al_c17b7119 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[7]));
  AL_DFF_X al_2d1290f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cbee0ff9[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da03ca6b[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_f508ac23 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[0]),
    .d(al_da03ca6b[1]),
    .e(al_da03ca6b[2]),
    .f(al_da03ca6b[3]),
    .o(al_a614d965));
  AL_MAP_LUT5 #(
    .EQN("((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(A)*~(E)+(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*~(E)+~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*A*E+(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*E)"),
    .INIT(32'haaaaf0cc))
    al_a3370975 (
    .a(al_4559aa8f),
    .b(al_a614d965),
    .c(al_4b0ede28),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_19b5d2a2[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff0ccaa00f0ccaa))
    al_950826ec (
    .a(al_7f73cd24),
    .b(al_da90d6e3),
    .c(al_3f457ae0),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .f(al_da03ca6b[22]),
    .o(al_19b5d2a2[10]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff0ccaa00f0ccaa))
    al_c602e9b9 (
    .a(al_695678a9),
    .b(al_9be05a01),
    .c(al_8f7d8418),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .f(al_da03ca6b[22]),
    .o(al_19b5d2a2[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7210a6f3 (
    .a(al_8a0179a4),
    .b(al_d7a13544),
    .c(al_b029b709[2]),
    .o(al_cbac66be));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_fffb8845 (
    .a(al_a6f911fa),
    .b(al_b029b709[2]),
    .c(al_da03ca6b[22]),
    .o(al_c4b36f25));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ee8b3376 (
    .a(al_cbac66be),
    .b(al_c4b36f25),
    .c(al_b029b709[3]),
    .o(al_19b5d2a2[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_5c6de1c3 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[13]),
    .d(al_da03ca6b[14]),
    .e(al_da03ca6b[15]),
    .f(al_da03ca6b[16]),
    .o(al_124b3a01));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_5b15f921 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[17]),
    .d(al_da03ca6b[18]),
    .e(al_da03ca6b[19]),
    .f(al_da03ca6b[20]),
    .o(al_b6c514a3));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d1c43482 (
    .a(al_124b3a01),
    .b(al_b6c514a3),
    .c(al_b029b709[2]),
    .o(al_a4ba3987));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D)*~((~C*~B*~A))+E*D*~((~C*~B*~A))+~(E)*D*(~C*~B*~A)+E*D*(~C*~B*~A))"),
    .INIT(32'hfffe0100))
    al_f2a8738d (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_b029b709[2]),
    .d(al_da03ca6b[21]),
    .e(al_da03ca6b[22]),
    .o(al_dacf88bd));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d1b0cfb3 (
    .a(al_a4ba3987),
    .b(al_dacf88bd),
    .c(al_b029b709[3]),
    .o(al_19b5d2a2[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_83c858 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[14]),
    .d(al_da03ca6b[15]),
    .e(al_da03ca6b[16]),
    .f(al_da03ca6b[17]),
    .o(al_da90d6e3));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_ff43f1f9 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[18]),
    .d(al_da03ca6b[19]),
    .e(al_da03ca6b[20]),
    .f(al_da03ca6b[21]),
    .o(al_3f457ae0));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(E)*~(D)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*~(D)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*E*D+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*D)"),
    .INIT(32'hffca00ca))
    al_f5e36baa (
    .a(al_da90d6e3),
    .b(al_3f457ae0),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .e(al_da03ca6b[22]),
    .o(al_19b5d2a2[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_f42ebbde (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[15]),
    .d(al_da03ca6b[16]),
    .e(al_da03ca6b[17]),
    .f(al_da03ca6b[18]),
    .o(al_9be05a01));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_8a07653e (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[19]),
    .d(al_da03ca6b[20]),
    .e(al_da03ca6b[21]),
    .f(al_da03ca6b[22]),
    .o(al_8f7d8418));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(E)*~(D)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*~(D)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*E*D+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*D)"),
    .INIT(32'hffca00ca))
    al_809ae8a7 (
    .a(al_9be05a01),
    .b(al_8f7d8418),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .e(al_da03ca6b[22]),
    .o(al_19b5d2a2[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_1d6fca89 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[16]),
    .d(al_da03ca6b[17]),
    .e(al_da03ca6b[18]),
    .f(al_da03ca6b[19]),
    .o(al_d7a13544));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    al_afcd213c (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[20]),
    .d(al_da03ca6b[21]),
    .e(al_da03ca6b[22]),
    .o(al_a6f911fa));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(E)*~(D)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*~(D)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*E*D+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*D)"),
    .INIT(32'hffca00ca))
    al_d54354c3 (
    .a(al_d7a13544),
    .b(al_a6f911fa),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .e(al_da03ca6b[22]),
    .o(al_19b5d2a2[16]));
  AL_MAP_LUT6 #(
    .EQN("(A*~((F*~(E)*~((~C*~B))+F*E*~((~C*~B))+~(F)*E*(~C*~B)+F*E*(~C*~B)))*~(D)+A*(F*~(E)*~((~C*~B))+F*E*~((~C*~B))+~(F)*E*(~C*~B)+F*E*(~C*~B))*~(D)+~(A)*(F*~(E)*~((~C*~B))+F*E*~((~C*~B))+~(F)*E*(~C*~B)+F*E*(~C*~B))*D+A*(F*~(E)*~((~C*~B))+F*E*~((~C*~B))+~(F)*E*(~C*~B)+F*E*(~C*~B))*D)"),
    .INIT(64'hffaafcaa03aa00aa))
    al_3d1c7ed1 (
    .a(al_b6c514a3),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_b029b709[2]),
    .e(al_da03ca6b[21]),
    .f(al_da03ca6b[22]),
    .o(al_60425dcb));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_6aa39fdd (
    .a(al_60425dcb),
    .b(al_b029b709[3]),
    .c(al_da03ca6b[22]),
    .o(al_19b5d2a2[17]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A)*~((~C*~B))+D*A*~((~C*~B))+~(D)*A*(~C*~B)+D*A*(~C*~B))"),
    .INIT(16'hfe02))
    al_f11425c4 (
    .a(al_3f457ae0),
    .b(al_b029b709[2]),
    .c(al_b029b709[3]),
    .d(al_da03ca6b[22]),
    .o(al_19b5d2a2[18]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A)*~((~C*~B))+D*A*~((~C*~B))+~(D)*A*(~C*~B)+D*A*(~C*~B))"),
    .INIT(16'hfe02))
    al_9cb67962 (
    .a(al_8f7d8418),
    .b(al_b029b709[2]),
    .c(al_b029b709[3]),
    .d(al_da03ca6b[22]),
    .o(al_19b5d2a2[19]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_d3306d47 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[1]),
    .d(al_da03ca6b[2]),
    .e(al_da03ca6b[3]),
    .f(al_da03ca6b[4]),
    .o(al_5976b207));
  AL_MAP_LUT5 #(
    .EQN("((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(A)*~(E)+(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*~(E)+~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*A*E+(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*E)"),
    .INIT(32'haaaaf0cc))
    al_63535bfb (
    .a(al_3a11d010),
    .b(al_5976b207),
    .c(al_1aa4ae3e),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_19b5d2a2[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_71d42eeb (
    .a(al_c4b36f25),
    .b(al_b029b709[3]),
    .c(al_da03ca6b[22]),
    .o(al_19b5d2a2[20]));
  AL_MAP_LUT6 #(
    .EQN("(F*~(E)*~((~D*~C*~B*~A))+F*E*~((~D*~C*~B*~A))+~(F)*E*(~D*~C*~B*~A)+F*E*(~D*~C*~B*~A))"),
    .INIT(64'hfffffffe00010000))
    al_33a4d6aa (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .e(al_da03ca6b[21]),
    .f(al_da03ca6b[22]),
    .o(al_19b5d2a2[21]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_1f275c9 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[2]),
    .d(al_da03ca6b[3]),
    .e(al_da03ca6b[4]),
    .f(al_da03ca6b[5]),
    .o(al_f5e8ffb7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccaaaaff000f0f))
    al_89375411 (
    .a(al_7f73cd24),
    .b(al_da90d6e3),
    .c(al_f5e8ffb7),
    .d(al_f35b497d),
    .e(al_b029b709[2]),
    .f(al_b029b709[3]),
    .o(al_19b5d2a2[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_5c9982ed (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[3]),
    .d(al_da03ca6b[4]),
    .e(al_da03ca6b[5]),
    .f(al_da03ca6b[6]),
    .o(al_66f5623c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccaaaaff000f0f))
    al_27466c83 (
    .a(al_695678a9),
    .b(al_9be05a01),
    .c(al_66f5623c),
    .d(al_b1cdfbfa),
    .e(al_b029b709[2]),
    .f(al_b029b709[3]),
    .o(al_19b5d2a2[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_c6706b40 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[4]),
    .d(al_da03ca6b[5]),
    .e(al_da03ca6b[6]),
    .f(al_da03ca6b[7]),
    .o(al_4b0ede28));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(E)+(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(E)+~((C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*E+(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*E)"),
    .INIT(32'haaaaccf0))
    al_f0b9382a (
    .a(al_cbac66be),
    .b(al_24ebd63f),
    .c(al_4b0ede28),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_19b5d2a2[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_1c07187a (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[5]),
    .d(al_da03ca6b[6]),
    .e(al_da03ca6b[7]),
    .f(al_da03ca6b[8]),
    .o(al_1aa4ae3e));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(E)+(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(E)+~((C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*E+(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*E)"),
    .INIT(32'haaaaccf0))
    al_480488b4 (
    .a(al_a4ba3987),
    .b(al_da6a2c78),
    .c(al_1aa4ae3e),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_19b5d2a2[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_9d5fdc6e (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[10]),
    .d(al_da03ca6b[11]),
    .e(al_da03ca6b[12]),
    .f(al_da03ca6b[13]),
    .o(al_7f73cd24));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_44bf2c04 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[6]),
    .d(al_da03ca6b[7]),
    .e(al_da03ca6b[8]),
    .f(al_da03ca6b[9]),
    .o(al_f35b497d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00ccccaaaaf0f0))
    al_5adb64b4 (
    .a(al_7f73cd24),
    .b(al_da90d6e3),
    .c(al_f35b497d),
    .d(al_3f457ae0),
    .e(al_b029b709[2]),
    .f(al_b029b709[3]),
    .o(al_19b5d2a2[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_2505f162 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[11]),
    .d(al_da03ca6b[12]),
    .e(al_da03ca6b[13]),
    .f(al_da03ca6b[14]),
    .o(al_695678a9));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_d5df933d (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[7]),
    .d(al_da03ca6b[8]),
    .e(al_da03ca6b[9]),
    .f(al_da03ca6b[10]),
    .o(al_b1cdfbfa));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00ccccaaaaf0f0))
    al_7a47b5f7 (
    .a(al_695678a9),
    .b(al_9be05a01),
    .c(al_b1cdfbfa),
    .d(al_8f7d8418),
    .e(al_b029b709[2]),
    .f(al_b029b709[3]),
    .o(al_19b5d2a2[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_5197f55 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[8]),
    .d(al_da03ca6b[9]),
    .e(al_da03ca6b[10]),
    .f(al_da03ca6b[11]),
    .o(al_24ebd63f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_1da461f7 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[12]),
    .d(al_da03ca6b[13]),
    .e(al_da03ca6b[14]),
    .f(al_da03ca6b[15]),
    .o(al_8a0179a4));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c9d81a24 (
    .a(al_24ebd63f),
    .b(al_8a0179a4),
    .c(al_b029b709[2]),
    .o(al_4559aa8f));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E)"),
    .INIT(32'hf0ccaaaa))
    al_73cf2530 (
    .a(al_4559aa8f),
    .b(al_d7a13544),
    .c(al_a6f911fa),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_19b5d2a2[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_f0f04691 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_da03ca6b[9]),
    .d(al_da03ca6b[10]),
    .e(al_da03ca6b[11]),
    .f(al_da03ca6b[12]),
    .o(al_da6a2c78));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f092bddc (
    .a(al_da6a2c78),
    .b(al_124b3a01),
    .c(al_b029b709[2]),
    .o(al_3a11d010));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_859ab835 (
    .a(al_3a11d010),
    .b(al_60425dcb),
    .c(al_b029b709[3]),
    .o(al_19b5d2a2[9]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    al_da111e4b (
    .a(al_4fb683a3),
    .b(al_36c58aac),
    .c(al_8c06569d),
    .d(num[0]),
    .o(al_c162c2a5));
  AL_DFF_X al_b353fbc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c162c2a5),
    .en(start),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3127e1e8));

endmodule 

