// Verilog netlist created by Tang Dynasty v5.6.71036
// Sat Oct 12 21:38:02 2024

`timescale 1ns / 1ps
module TEMAC_CORE
  (
  gmii_col,
  gmii_crs,
  gmii_rx_er,
  gmii_rx_vld,
  gmii_rxd,
  gmii_tx_clken,
  mac_cfg_vector,
  mdio_in,
  pause_req,
  pause_source_addr,
  pause_val,
  reset,
  rx_clk_en,
  rx_mac_clk,
  s_axi_aclk,
  s_axi_araddr,
  s_axi_arvalid,
  s_axi_awaddr,
  s_axi_awvalid,
  s_axi_bready,
  s_axi_rready,
  s_axi_wdata,
  s_axi_wvalid,
  tx_clk_en,
  tx_data,
  tx_data_en,
  tx_ifg_val,
  tx_mac_clk,
  tx_stop,
  unicast_addr,
  gmii_tx_en,
  gmii_tx_er,
  gmii_txd,
  mdio_clk,
  mdio_oen,
  mdio_out,
  rx_correct_frame,
  rx_data,
  rx_data_vld,
  rx_error_frame,
  rx_status_vector,
  rx_status_vld,
  s_axi_arready,
  s_axi_awready,
  s_axi_bresp,
  s_axi_bvalid,
  s_axi_rdata,
  s_axi_rresp,
  s_axi_rvalid,
  s_axi_wready,
  speed_10,
  speed_100,
  speed_1000,
  tx_collision,
  tx_rdy,
  tx_retransmit,
  tx_status_vector,
  tx_status_vld
  );

  input gmii_col;
  input gmii_crs;
  input gmii_rx_er;
  input gmii_rx_vld;
  input [7:0] gmii_rxd;
  input gmii_tx_clken;
  input [19:0] mac_cfg_vector;
  input mdio_in;
  input pause_req;
  input [47:0] pause_source_addr;
  input [15:0] pause_val;
  input reset;
  input rx_clk_en;
  input rx_mac_clk;
  input s_axi_aclk;
  input [7:0] s_axi_araddr;
  input s_axi_arvalid;
  input [7:0] s_axi_awaddr;
  input s_axi_awvalid;
  input s_axi_bready;
  input s_axi_rready;
  input [31:0] s_axi_wdata;
  input s_axi_wvalid;
  input tx_clk_en;
  input [7:0] tx_data;
  input tx_data_en;
  input [7:0] tx_ifg_val;
  input tx_mac_clk;
  input tx_stop;
  input [47:0] unicast_addr;
  output gmii_tx_en;
  output gmii_tx_er;
  output [7:0] gmii_txd;
  output mdio_clk;
  output mdio_oen;
  output mdio_out;
  output rx_correct_frame;
  output [7:0] rx_data;
  output rx_data_vld;
  output rx_error_frame;
  output [26:0] rx_status_vector;
  output rx_status_vld;
  output s_axi_arready;
  output s_axi_awready;
  output [1:0] s_axi_bresp;
  output s_axi_bvalid;
  output [31:0] s_axi_rdata;
  output [1:0] s_axi_rresp;
  output s_axi_rvalid;
  output s_axi_wready;
  output speed_10;
  output speed_100;
  output speed_1000;
  output tx_collision;
  output tx_rdy;
  output tx_retransmit;
  output [28:0] tx_status_vector;
  output tx_status_vld;

  parameter P_ADD_FILT_EN = 1'b1;
  parameter P_ADD_FILT_LIST = 3;
  parameter P_HALF_DUPLEX = 1'b1;
  parameter P_HOST_EN = 1'b1;
  parameter P_SPEED_1000 = 1'b0;
  parameter P_SPEED_10_100 = 1'b0;
  parameter P_TRI_SPEED = 1'b1;
  // localparam P_CLK_EN = 1'b1;
  wire [7:0] al_aeb75558;
  wire [4:0] al_47e69606;
  wire [4:0] al_2b21b090;
  wire [4:0] al_a6a28e17;
  wire [7:0] al_f6e00c9;
  wire [15:0] al_e1f88382;
  wire [15:0] al_e6e0b636;
  wire [15:0] al_7d74a9c;
  wire [7:0] al_9c49a375;
  wire [7:0] al_de1356f0;
  wire [4:0] al_67a4bdfd;
  wire [4:0] al_cade1083;
  wire [47:0] al_c5235ca5;
  wire [15:0] al_522cbac;
  wire [2:0] al_520772a3;
  wire  al_de41ced;
  wire  al_76834e7a;
  wire  al_bf066204;
  wire  al_84a2caa3;
  wire  al_cba22e49;
  wire [7:0] al_c01774ad;
  wire [15:0] al_64a46519;
  wire [15:0] al_f69b891;
  wire [15:0] al_8a4cc919;
  wire [5:0] al_a9476246;
  wire [5:0] al_81fd75dc;
  wire [14:0] al_5c90f2da;
  wire [7:0] al_eb34b0be;
  wire [3:0] al_6ae08f56;
  wire [3:0] al_f0ba390f;
  wire [3:0] al_2fda9ea8;
  wire [7:0] al_42702950;
  wire [7:0] al_3b8f6a2b;
  wire [11:0] al_302d0d8b;
  wire [3:0] al_ecabfff7;
  wire [3:0] al_18a8d68c;
  wire [3:0] al_e08d2b14;
  wire [3:0] al_2ddf456e;
  wire [3:0] al_55d8b8f7;
  wire [3:0] al_4c8ab20f;
  wire [3:0] al_e7fcc128;
  wire [7:0] al_f279ca9c;
  wire [7:0] al_be455f81;
  wire [7:0] al_53486c5d;
  wire [5:0] al_a60f8a1f;
  wire [5:0] al_c364719f;
  wire [7:0] al_eb5eeaf9;
  wire [7:0] al_6f6e3b4e;
  wire [7:0] al_60c7c349;
  wire [7:0] al_dbc70e2f;
  wire [31:0] al_fa4d6e00;
  wire [31:0] al_871e6587;
  wire [6:0] al_3f753490;
  wire [31:0] al_7de51101;
  wire [31:0] al_3cae1837;
  wire [31:0] al_4197a0a2;
  wire [31:0] al_42381c95;
  wire [31:0] al_ae69e57d;
  wire [31:0] al_a3c2ad2a;
  wire [31:0] al_1062ede0;
  wire [31:0] al_677d00f0;
  wire [31:0] al_9e3bc263;
  wire [31:0] al_e340ee08;
  wire [31:0] al_a100d2c5;
  wire [31:0] al_52b0078;
  wire [1:0] al_44560df6;
  wire [31:0] al_32c99495;
  wire [15:0] al_1cb63986;
  wire [5:0] al_71b90bfa;
  wire [15:0] al_81b839ee;
  wire [15:0] al_469f2a04;
  wire [15:0] al_ff43a01c;
  wire [7:0] al_1a0f7d2b;
  wire [31:0] al_53a2c384;
  wire [23:0] al_5f1c4763;
  wire [31:0] al_e57de54;
  wire [9:0] al_e023302;
  wire [9:0] al_7b9b882d;
  wire [9:0] al_5c2983f8;
  wire [15:0] al_1e120105;
  wire [15:0] al_ea827a0c;
  wire [15:0] al_4f3b20c;
  wire [14:0] al_b9d3b2c1;
  wire [14:0] al_9e843f7;
  wire [14:0] al_66bdfa10;
  wire [15:0] al_2814a16d;
  wire [15:0] al_13349257;
  wire [13:0] al_26b248e8;
  wire [1:0] al_b449eeb9;
  wire [7:0] al_583c216b;
  wire [7:0] al_1d03242c;
  wire [7:0] al_5e036bbd;
  wire [5:0] al_ef7f6f7b;
  wire [3:0] al_6aa6d3c8;
  wire [1:0] al_4ceb8d18;
  wire [24:0] al_36654522;
  wire [1:0] al_54280ae3;
  wire [15:0] al_ddf438c2;
  wire [15:0] al_6133949d;
  wire [15:0] al_bd413a73;
  wire [15:0] al_e799d30a;
  wire [15:0] al_33bfe5eb;
  wire [15:0] al_dd83fb37;
  wire [15:0] al_7bd9ce9a;
  wire [15:0] al_4c32576a;
  wire [9:0] al_aa981a62;
  wire [3:0] al_21330e1d;
  wire [14:0] al_90205973;
  wire [13:0] al_69384d3c;
  wire [3:0] al_a21ad81c;
  wire [3:0] al_acfeaf96;
  wire [4:0] al_64a47488;
  wire [2:0] al_fff0fd72;
  wire [2:0] al_471dc00c;
  wire [12:0] al_278aa6ae;
  wire [12:0] al_23bcf331;
  wire [13:0] al_56ef451f;
  wire [1:0] al_d2dd6034;
  wire [1:0] al_fd60fee0;
  wire [7:0] al_4228c99a;
  wire [5:0] al_c9168fb8;
  wire [5:0] al_55a9d56d;
  wire [3:0] al_30c5253d;
  wire [18:0] al_332a045d;
  wire [18:0] al_dbdaab6;
  wire [19:0] al_cc156ef4;
  wire [9:0] al_ab37059b;
  wire [14:0] al_618d6d02;
  wire [14:0] al_17c3d18e;
  wire [14:0] al_e29488b2;
  wire [14:0] al_1a83737a;
  wire [31:0] al_d62b96ee;
  wire [23:0] al_2be5d117;
  wire [31:0] al_e66356bf;
  wire [1:0] al_321109d3;
  wire [1:0] al_aea1aa30;
  wire [7:0] al_2ea27c82;
  wire [7:0] al_f5fe9553;
  wire [7:0] al_d275691c;
  wire [7:0] al_8b969422;
  wire [7:0] al_31841a5b;
  wire [7:0] al_da791a9b;
  wire [7:0] al_d567b233;
  wire [7:0] al_47ab7609;
  wire [7:0] al_2453f186;
  wire [7:0] al_d1fcb50b;
  wire [7:0] al_f24f9b58;
  wire [14:0] al_59a6ee8e;
  wire [14:0] al_49200bab;
  wire [15:0] al_83a6bf62;
  wire [10:0] al_1b8c3389;
  wire [10:0] al_ee979a13;
  wire [14:0] al_5305cb61;
  wire [14:0] al_b084da19;
  wire [14:0] al_b7d1cff2;
  wire [14:0] al_e31e36f5;
  wire [4:0] al_df9b9d5b;
  wire [7:0] al_18d64456;
  wire [7:0] al_5743d58d;
  wire [7:0] al_b2d09c6f;
  wire [13:0] al_1d28bc9;
  wire [7:0] al_6a6d2547;
  wire [7:0] al_3ac23457;
  wire [7:0] al_2e49f5b3;
  wire [3:0] al_1fc5093b;
  wire [1:0] al_3ab98f26;
  wire [1:0] al_9bde74c4;
  wire [9:0] al_3ce55a07;
  wire [9:0] al_2e44f12e;
  wire [9:0] al_302a167b;
  wire [15:0] al_eb2b30c3;
  wire [13:0] al_cb8cffb4;
  wire [2:0] al_2a1554ab;
  wire [2:0] al_cf2a0a44;
  wire [1:0] al_931288d8;
  wire [63:0] al_5ffd8cb3;
  wire [63:0] al_b7012aee;
  wire [63:0] al_f07b9ef6;
  wire [3:0] al_f931229;
  wire [31:0] al_4248a527;
  wire [2:0] al_7f29f8c;
  wire [2:0] al_abfa408b;
  wire [15:0] al_6a2b89f7;
  wire [127:0] al_d7778ec8;
  wire  al_aa714f0f;
  wire  al_50654b35;
  wire  al_554dd8ee;
  wire  al_51ce9e18;
  wire  al_5f7aacbd;
  wire  al_338c309a;
  wire  al_8345e39d;
  wire  al_d55c6f72;
  wire  al_37adc87c;
  wire  al_82d0eff2;
  wire  al_c6b2b040;
  wire  al_9a8f38a1;
  wire  al_86319e2;
  wire  al_b7ea58da;
  wire  al_b723aa66;
  wire  al_ae9f73b7;
  wire  al_5039df42;
  wire  al_40ffa4c8;
  wire  al_e739923;
  wire  al_62f30b7f;
  wire  al_11c347b2;
  wire  al_c4aea171;
  wire  al_4753a8f9;
  wire  al_68f10ad3;
  wire  al_38bca4e9;
  wire  al_a1ae1d55;
  wire  al_8272529a;
  wire  al_7bcaf633;
  wire  al_c0e589a5;
  wire  al_ffaac04;
  wire  al_f510713e;
  wire  al_44266b04;
  wire  al_c183d3b1;
  wire  al_5d766886;
  wire  al_743eaea9;
  wire  al_429251b;
  wire  al_39cac231;
  wire  al_8f559a59;
  wire  al_53e610e6;
  wire  al_c246767f;
  wire  al_a5ba552b;
  wire  al_6b621a04;
  wire  al_d2549f15;
  wire  al_5a10d00d;
  wire  al_9fedaeeb;
  wire  al_f1b5d549;
  wire  al_803791d8;
  wire  al_e06bf58f;
  wire  al_6ce7e86b;
  wire  al_f75db11b;
  wire  al_f46dd33d;
  wire  al_899c7875;
  wire  al_9ca6a99d;
  wire  al_83bf8364;
  wire  al_25b9d53e;
  wire  al_66f1c0a9;
  wire  al_95b2c02e;
  wire  al_df1c692d;
  wire  al_f951c654;
  wire [47:0] al_b091d0de;
  wire [47:0] al_e49fcd23;
  wire  al_f0b71806;
  wire  al_593a2319;
  wire  al_8dea866b;
  wire  al_f5169e61;
  wire  al_ee3af5c0;
  wire  al_928a2d4f;
  wire  al_5995850b;
  wire  al_70bede4a;
  wire  al_58cfbf60;
  wire  al_fe6f17e2;
  wire  al_11243436;
  wire  al_b7c18d6c;
  wire  al_f383744d;
  wire  al_8dce46fa;
  wire  al_85cd42a7;
  wire  al_3e863ba;
  wire  al_2c55a3d3;
  wire  al_e4cf91e2;
  wire  al_5d5dee64;
  wire  al_7ff105dd;
  wire  al_c32e7d0;
  wire  al_e6a1e4d5;
  wire  al_e2546db0;
  wire  al_33bf9b84;
  wire  al_aa8be9ce;
  wire  al_9f180be0;
  wire  al_7c64c6fa;
  wire  al_cafe8108;
  wire  al_cd2ca50c;
  wire  al_b28e21a8;
  wire  al_2379dade;
  wire  al_13b54967;
  wire [7:0] al_e8711ae2;
  wire [47:0] al_9207c009;
  wire [47:0] al_ddb70824;
  wire [47:0] al_f1ef691c;
  wire [47:0] al_1c1c7167;
  wire al_bd973c28;
  wire al_a9188fac;
  wire al_29be6517;
  wire al_31b957f1;
  wire al_2dd67b98;
  wire al_816cf877;
  wire al_a69b9244;
  wire al_ce6f4d2;
  wire al_8868df5f;
  wire al_54d1791f;
  wire al_2e24cdc2;
  wire al_40609b11;
  wire al_67528d08;
  wire al_75607bc2;
  wire al_bcfe99bb;
  wire al_82b20445;
  wire al_c7af49f0;
  wire al_3bed0c06;
  wire al_43bc4712;
  wire al_6b1e934b;
  wire al_43f140b9;
  wire al_f5fab0c0;
  wire al_613f9025;
  wire al_9149a8cc;
  wire al_502a557a;
  wire al_f84368bb;
  wire al_a57398e0;
  wire al_cad59eac;
  wire al_157db10;
  wire al_b6be6226;
  wire al_fb677f9;
  wire al_12adcf0d;
  wire al_9d0e1a05;
  wire al_12c00371;
  wire al_1cb53946;
  wire al_414fb589;
  wire al_8bc3cc10;
  wire al_8ae11e67;
  wire al_5ea7feee;
  wire al_b4de44d1;
  wire al_c00b14c1;
  wire al_67c63555;
  wire al_f655e852;
  wire al_2086e64;
  wire al_cad879da;
  wire al_51967b89;
  wire al_fe18e71f;
  wire al_aad3b572;
  wire al_14a7b701;
  wire al_f41510c0;
  wire al_74fb81be;
  wire al_1f397d18;
  wire al_b7dabd2c;
  wire al_d0814789;
  wire al_5686da25;
  wire al_58fac850;
  wire al_732c5a74;
  wire al_e545d06c;
  wire al_93727b8b;
  wire al_1ca59da3;
  wire al_6c3542a2;
  wire al_b0dc2f75;
  wire al_389c7bee;
  wire al_98c25345;
  wire al_bd3e169c;
  wire al_b821ca29;
  wire al_16302c3d;
  wire al_60057698;
  wire al_44dddc1d;
  wire al_d32c67d0;
  wire al_31529785;
  wire al_e48259f9;
  wire al_7b681f71;
  wire al_51616140;
  wire al_c9465832;
  wire al_5b289734;
  wire al_c2520419;
  wire al_f164e0a;
  wire al_74354c6e;
  wire al_c292362f;
  wire al_5b37fe28;
  wire al_e101ff9a;
  wire al_aaead9c7;
  wire al_a6ff135b;
  wire al_5a6020b4;
  wire al_82120dcc;
  wire al_4dabd984;
  wire al_430719be;
  wire al_e18e0a15;
  wire al_2de0dbf6;
  wire al_c2be7784;
  wire al_a523c2cb;
  wire al_b2deb19c;
  wire al_6bdd801e;
  wire al_b2b271cb;
  wire al_4d9c2a7a;
  wire al_18e5b9af;
  wire al_93abd71;
  wire al_3a74e04b;
  wire al_33e46ce3;
  wire al_47f8fdc1;
  wire al_6b96fb99;
  wire al_f55c93aa;
  wire al_1bba34ee;
  wire al_82835dec;
  wire al_eb74cd21;
  wire al_fb8448e4;
  wire al_e2a1fab3;
  wire al_511fc342;
  wire al_7f616b69;
  wire al_c192e229;
  wire al_5ecede8f;
  wire al_90044ea4;
  wire al_4b956df0;
  wire al_a88739b8;
  wire al_eeb871e3;
  wire al_b93d302f;
  wire al_fd543856;
  wire al_abceb3af;
  wire al_d9c2bbe5;
  wire al_1a69e04c;
  wire al_4940717b;
  wire al_65719225;
  wire al_5d511a0d;
  wire al_1da67580;
  wire al_889a47a2;
  wire al_b306469e;
  wire al_6aba2287;
  wire al_7fd108f9;
  wire al_a51041a6;
  wire al_d78ef14f;
  wire al_5097d6f;
  wire al_b65ba3d5;
  wire al_9eb158b7;
  wire al_1421d0c8;
  wire al_d7389040;
  wire al_ac2b4841;
  wire al_69e62d6a;
  wire al_5e18973f;
  wire al_fe501ed1;
  wire al_d1c7d2fd;
  wire al_95c95cdd;
  wire al_7dd23876;
  wire al_b3b32038;
  wire al_a655b507;
  wire al_758baf6a;
  wire al_f4206233;
  wire al_82c4c889;
  wire al_1c26630b;
  wire al_38ceef8c;
  wire al_7c925305;
  wire al_41a3eebf;
  wire al_5b5454d7;
  wire al_a52c4218;
  wire al_2456cab6;
  wire al_c88ff5bc;
  wire al_d7c1f764;
  wire al_ca164e15;
  wire al_6fc51898;
  wire al_460e3807;
  wire al_b1302323;
  wire al_2f1e9be;
  wire al_5617038b;
  wire al_7807b4dd;
  wire al_511c2516;
  wire al_c4a95f07;
  wire al_452dacc5;
  wire al_9cae7666;
  wire al_495ac57d;
  wire al_d811a788;
  wire al_8e5a365f;
  wire al_2c74b50c;
  wire al_c92c521a;
  wire al_f9514cde;
  wire al_da725511;
  wire al_23e59594;
  wire al_d133c6bf;
  wire al_de6e30a1;
  wire al_fbe1feab;
  wire al_240f6a60;
  wire al_58e61c93;
  wire al_6127633d;
  wire al_a7dbaac0;
  wire al_e495ee45;
  wire al_16d49820;
  wire al_a76fca28;
  wire al_f2e8c346;
  wire al_715e8e22;
  wire al_5a4539df;
  wire al_637ddda1;
  wire al_d811499f;
  wire al_53653f1d;
  wire al_9848ae60;
  wire al_d19ca65b;
  wire al_aceaab6b;
  wire al_e78cfe9;
  wire al_d5fb3fbb;
  wire al_18862d32;
  wire al_fb84638b;
  wire al_78920a9b;
  wire al_6298ef12;
  wire al_38ea65b9;
  wire al_124a5ff1;
  wire al_6842e259;
  wire al_524c4c86;
  wire al_2d0b2d41;
  wire al_7ca091b;
  wire al_e1e36fb;
  wire al_f4745b25;
  wire al_a533f139;
  wire al_38a4dea8;
  wire al_2839f3fc;
  wire al_16bdb356;
  wire al_1b4e1994;
  wire al_a2b6b866;
  wire al_8f160d47;
  wire al_a0ae817c;
  wire al_f6f1aa20;
  wire al_b436d586;
  wire al_197bd181;
  wire al_10c967cd;
  wire al_df75d779;
  wire al_587464d;
  wire al_fec67178;
  wire al_713dc35e;
  wire al_22f0d00f;
  wire al_33156af5;
  wire al_8f006d4e;
  wire al_de5e814a;
  wire al_eb5ace4a;
  wire al_902ad644;
  wire al_c5eafaca;
  wire al_63772beb;
  wire al_69a4217a;
  wire al_525bf098;
  wire al_f55cb982;
  wire al_d1b2b221;
  wire al_aa6b82f0;
  wire al_66d7ef91;
  wire al_4462abf6;
  wire al_ca7097d4;
  wire al_48f0356f;
  wire al_e9410de9;
  wire al_90130b74;
  wire al_30591f5d;
  wire al_760b1195;
  wire al_22e99ffa;
  wire al_b936a4eb;
  wire al_16296d60;
  wire al_fb466fd8;
  wire al_6fbcf05d;
  wire al_c5d247c0;
  wire al_b3b873e8;
  wire al_5d24a167;
  wire al_d4b6c586;
  wire al_240a1ace;
  wire al_27fc47ee;
  wire al_d38bd427;
  wire al_ffb977ef;
  wire al_c7821d7e;
  wire al_ec112ad9;
  wire al_1ff3d4e5;
  wire al_68cc6b50;
  wire al_d7515c44;
  wire al_39b879bd;
  wire al_dd95f235;
  wire al_41fb49d4;
  wire al_937f8e6e;
  wire al_d1b5a8f4;
  wire al_f6f8b1fe;
  wire al_fcdf9700;
  wire al_919f4410;
  wire al_8a13cd79;
  wire al_38bb9e5e;
  wire al_efdfec25;
  wire al_a2d51717;
  wire al_594ca757;
  wire al_e2aa4ae4;
  wire al_f4b9a391;
  wire al_8b7519f2;
  wire al_1883a4da;
  wire al_f947ca8;
  wire al_60adcd8c;
  wire al_618a5a5f;
  wire al_1c6af38a;
  wire al_b3550f8b;
  wire al_852e5bbe;
  wire al_ee5f9e50;
  wire al_a1c88bcd;
  wire al_4a8487b2;
  wire al_72a9a166;
  wire al_b58b5a6;
  wire al_6cc2d7f5;
  wire al_71411c23;
  wire al_56e2186e;
  wire al_9e23e23c;
  wire al_f423313d;
  wire al_ef0c62ea;
  wire al_46dd4bfb;
  wire al_4db0ca34;
  wire al_39575073;
  wire al_5ecd0d98;
  wire al_b809a0d;
  wire al_488ce459;
  wire al_2acb5425;
  wire al_8e73257f;
  wire al_36260f8d;
  wire al_1d55dde3;
  wire al_66a27b74;
  wire al_69ac11ac;
  wire al_bdab8dd4;
  wire al_2156b30e;
  wire al_55bc11eb;
  wire al_665205be;
  wire al_450a8cba;
  wire al_b14c08d7;
  wire al_14c1bc93;
  wire al_9cc4302;
  wire al_31ede2e2;
  wire al_c291f47d;
  wire al_b37ae739;
  wire al_b8f3be80;
  wire al_cee59967;
  wire al_8ba03385;
  wire al_9ec235f9;
  wire al_76f4f274;
  wire al_8b9cbde3;
  wire al_4ebb1964;
  wire al_a4aaca2e;
  wire al_b93f6564;
  wire al_655c284a;
  wire al_e1f066de;
  wire al_5a17606d;
  wire al_26874532;
  wire al_a360ff8;
  wire al_7fda1410;
  wire al_4f925611;
  wire al_7f161bf2;
  wire al_9d802914;
  wire al_830d7e;
  wire al_27f7f6ec;
  wire al_afd5fd5d;
  wire al_6a277bd4;
  wire al_f1c0fe91;
  wire al_18128b53;
  wire al_12c9315c;
  wire al_54829ae8;
  wire al_7360a7c0;
  wire al_5cbbf9cd;
  wire al_2d86aa6e;
  wire al_63df2227;
  wire al_12b617e9;
  wire al_77c268d4;
  wire al_aecc1a53;
  wire al_46fb2129;
  wire al_6492ae8;
  wire al_9e9040d4;
  wire al_f44ba8da;
  wire al_adf2eefc;
  wire al_944f1baf;
  wire al_ee5a9fb;
  wire al_15e31402;
  wire al_955255ce;
  wire al_61af39ad;
  wire al_20afe6c0;
  wire al_138eaec3;
  wire al_72045a1c;
  wire al_ee917930;
  wire al_88c12a03;
  wire al_ddac5e8d;
  wire al_5d42041c;
  wire al_f78634c8;
  wire al_33d9db52;
  wire al_6b647f54;
  wire al_c3ba6eaa;
  wire al_338b9100;
  wire al_fabf91f7;
  wire al_2169fa2d;
  wire al_a698f8f;
  wire al_14067aef;
  wire al_c0936433;
  wire al_86bf0006;
  wire al_8bef06bd;
  wire al_27629aac;
  wire al_3560f04f;
  wire al_ae3e538d;
  wire al_a15918b4;
  wire al_60f51d47;
  wire al_9439ddc;
  wire al_b3220547;
  wire al_b8f86eed;
  wire al_b0b9c021;
  wire al_8cebb59e;
  wire al_4ab032f9;
  wire al_72bd37a4;
  wire al_b2e646bb;
  wire al_18642257;
  wire al_a37dea2d;
  wire al_41d2ce29;
  wire al_e5a67968;
  wire al_39c05299;
  wire al_dd43c64f;
  wire al_1bdd94f8;
  wire al_8f689368;
  wire al_d6baa558;
  wire al_7ac96e46;
  wire al_9a2dcc24;
  wire al_4c9b2533;
  wire al_c5450b82;
  wire al_4696ac48;
  wire al_7710deab;
  wire al_e1057698;
  wire al_d6bd6336;
  wire al_c99d4c23;
  wire al_82dda9be;
  wire al_9cabf6c6;
  wire al_225d06ad;
  wire al_74c05d28;
  wire al_1ce99d34;
  wire al_6c6d3d88;
  wire al_597cc1f6;
  wire al_d83e61fb;
  wire al_932a07c7;
  wire al_7ffbbf6e;
  wire al_7a7628f9;
  wire al_ebdfe328;
  wire al_7c1aee64;
  wire al_cb67e17c;
  wire al_5274ea30;
  wire al_4e1502ae;
  wire al_48908c7b;
  wire al_cc7e79c9;
  wire al_91fb7c78;
  wire al_e646046;
  wire al_3ccf053a;
  wire al_5107a44a;
  wire al_4409fb45;
  wire al_b605ded6;
  wire al_b70fe470;
  wire al_124e348a;
  wire al_d671f8ef;
  wire al_e34977fd;
  wire al_c611b356;
  wire al_e890f462;
  wire al_b610aa54;
  wire al_a3a88d3f;
  wire al_f00de1fc;
  wire al_d9299255;
  wire al_88bee87;
  wire al_c57a154;
  wire al_32ab2441;
  wire al_9613edfd;
  wire al_d7a47bf6;
  wire al_8b0ea091;
  wire al_f0d27177;
  wire al_ce4327dc;
  wire al_13cf5eba;
  wire al_46839cba;
  wire al_bbbfb344;
  wire al_66f2b6b8;
  wire al_2eea7a5a;
  wire al_f3170c9;
  wire al_2270269f;
  wire al_179ef786;
  wire al_df30c316;
  wire al_ba6d5331;
  wire al_1fad8912;
  wire al_38e61a96;
  wire al_43d0de98;
  wire al_36b29f2;
  wire al_d4a11187;
  wire al_12dfe9dc;
  wire al_75def4ef;
  wire al_aa9f8872;
  wire al_153d6f9e;
  wire al_44348d99;
  wire al_134f4cf5;
  wire al_21b2c715;
  wire al_6f75ef0e;
  wire al_b95885c7;
  wire al_49b1129;
  wire al_decf41ac;
  wire al_d49fbba9;
  wire al_c4d37b2;
  wire al_1dcf5c5b;
  wire al_45a6c91;
  wire al_7c20ee3b;
  wire al_2ac16c9f;
  wire al_f5080327;
  wire al_e9f83d6e;
  wire al_81378cfb;
  wire al_31415f80;
  wire al_3f4108ac;
  wire al_f02638e3;
  wire al_60b3be17;
  wire al_25af80c5;
  wire al_96064004;
  wire al_f9a0f4e;
  wire al_95894036;
  wire al_6fed1e72;
  wire al_8f867af4;
  wire al_f03499fc;
  wire al_db3e7a3b;
  wire al_f1799bbf;
  wire al_c5cae25a;
  wire al_6f517dcb;
  wire al_5d55f7bd;
  wire al_93f12ca5;
  wire al_822d50d7;
  wire al_be626253;
  wire al_55aaf816;
  wire al_a5f70472;
  wire al_5c2a2da8;
  wire al_65f65cdd;
  wire al_6b3de12e;
  wire al_30e55692;
  wire al_efa05a0c;
  wire al_1e582b4d;
  wire al_9c659f6;
  wire al_3e9eebf5;
  wire al_384019b7;
  wire al_abdbe49;
  wire al_b3d5e449;
  wire al_5c7d4b11;
  wire al_a468a88f;
  wire al_ae1bb7ab;
  wire al_ba174b4c;
  wire al_fdc321a5;
  wire al_bc9d849e;
  wire al_42c40cf0;
  wire al_a095939;
  wire al_8a98fa0e;
  wire al_df322506;
  wire al_9a3d38d8;
  wire al_ac4196c0;
  wire al_dacf8588;
  wire al_509509ae;
  wire al_13154bf6;
  wire al_e1dab4c9;
  wire al_336d8f19;
  wire al_9f21cd24;
  wire al_b242277f;
  wire al_16c52309;
  wire al_ec602117;
  wire al_162f415f;
  wire al_c862ea52;
  wire al_f9e26d2b;
  wire al_d1bf4e26;
  wire al_adf11663;
  wire al_b8530805;
  wire al_3fdafe26;
  wire al_ff7075f1;
  wire al_1b7fc148;
  wire al_109f9c2b;
  wire al_c758ee36;
  wire al_8c3b9f16;
  wire al_ea736991;
  wire al_31cc16da;
  wire al_29cb9079;
  wire al_6f2b16fe;
  wire al_46118f46;
  wire al_f97fd11e;
  wire al_4c3c2401;
  wire al_a409c88e;
  wire al_4360005c;
  wire al_e2dc2eea;
  wire al_f0362cc;
  wire al_4f800f89;
  wire al_d5a6be8d;
  wire al_4d5dd241;
  wire al_ce94a07b;
  wire al_6598ce3a;
  wire al_9e79b57b;
  wire al_2c3ff84c;
  wire al_b1f059e9;
  wire al_5d14a06f;
  wire al_debb55eb;
  wire al_9b66e5cd;
  wire al_e729b3e2;
  wire al_9f6030e;
  wire al_b9b188f3;
  wire al_8fc9814c;
  wire al_b99dff45;
  wire al_50559550;
  wire al_6e672ebc;
  wire al_b19043fc;
  wire al_fd106601;
  wire al_ca4883db;
  wire al_db678397;
  wire al_cb7ab50c;
  wire al_9809ce8b;
  wire al_62730356;
  wire al_5b221454;
  wire al_53cf6c8d;
  wire al_72818778;
  wire al_7d123240;
  wire al_58a58247;
  wire al_379fd30a;
  wire al_fea77e50;
  wire al_156e79c6;
  wire al_9fbc578a;
  wire al_ceee241e;
  wire al_a71f4bd6;
  wire al_a296c440;
  wire al_2dbca608;
  wire al_aff8bba6;
  wire al_73bb0740;
  wire al_a231fc3f;
  wire al_9ff01b51;
  wire al_4e287126;
  wire al_5e767b18;
  wire al_46f6a926;
  wire al_1ea4ba5b;
  wire al_de9cd38;
  wire al_b1d9ebd5;
  wire al_b0d5abbb;
  wire al_95293982;
  wire al_9ac9e635;
  wire al_e7bc5d6e;
  wire al_c68f2ca9;
  wire al_81a5ac08;
  wire al_d424a202;
  wire al_aaec830f;
  wire al_7680e48;
  wire al_cb6844a5;
  wire al_b53d4bb7;
  wire al_1093568b;
  wire al_720c32ab;
  wire al_cd4fb40c;
  wire al_174be6c3;
  wire al_24bcb54c;
  wire al_35d72057;
  wire al_ef9c2399;
  wire al_17a2b8b;
  wire al_da621072;
  wire al_7680352d;
  wire al_c5272fc1;
  wire al_ff9a0466;
  wire al_3cb62398;
  wire al_ba6a9a7d;
  wire al_459462b6;
  wire al_143a100;
  wire al_8ce032ae;
  wire al_e7ec627;
  wire al_d8e2b166;
  wire al_f2be847d;
  wire al_8eaf8008;
  wire al_22412e0c;
  wire al_4210af67;
  wire al_2be5cde7;
  wire al_279abee0;
  wire al_b8bd8e77;
  wire al_1f78cc6;
  wire al_b42ee6d4;
  wire al_856accff;
  wire al_4952d975;
  wire al_86ce862e;
  wire al_d5178990;
  wire al_9a990f97;
  wire al_a7784e58;
  wire al_3009e595;
  wire al_c75b827e;
  wire al_968a4ecb;
  wire al_26e81f34;
  wire al_9ea76e6c;
  wire al_63060b04;
  wire al_3171227d;
  wire al_360de72;
  wire al_e707cc0b;
  wire al_84db4232;
  wire al_6a7aee90;
  wire al_af35a257;
  wire al_7fda34f5;
  wire al_318f23df;
  wire al_8202a39;
  wire al_33069608;
  wire al_b430139c;
  wire al_5ce3a1c4;
  wire al_e7b257ab;
  wire al_8a331b5c;
  wire al_221dcc8d;
  wire al_396e35f3;
  wire al_c34e4fd4;
  wire al_57958b12;
  wire al_3d6f4ec0;
  wire al_7dd043ee;
  wire al_3226aea6;
  wire al_54e1a5bd;
  wire al_9d8455d9;
  wire al_7a415511;
  wire al_26f9894f;
  wire al_ef281c2d;
  wire al_1db814d4;
  wire al_525a0f14;
  wire al_3829c8d6;
  wire al_c5560662;
  wire al_26c32275;
  wire al_df53a2ee;
  wire al_a0dade4c;
  wire al_eb84a31d;
  wire al_fe26d7bb;
  wire al_7a228cbe;
  wire al_be8ce4c3;
  wire al_bdda766f;
  wire al_16346f67;
  wire al_90aba52e;
  wire al_b4b4f932;
  wire al_39bec123;
  wire al_6819cc15;
  wire al_22cdf2f;
  wire al_1c995ac6;
  wire al_2ef83128;
  wire al_2cadd0ad;
  wire al_facb0130;
  wire al_3bd7786d;
  wire al_f32db70e;
  wire al_d4f4862c;
  wire al_d991794b;
  wire al_78564a3b;
  wire al_f3a13de0;
  wire al_b06018b7;
  wire al_537f614b;
  wire al_c89ba6ec;
  wire al_19aaf769;
  wire al_35dbcd92;
  wire al_6a936812;
  wire al_cc204c06;
  wire al_f5e85a1;
  wire al_1520e86d;
  wire al_47214dbf;
  wire al_5c754024;
  wire al_8e143433;
  wire al_3e1806d9;
  wire al_567c0900;
  wire al_ee8c5e52;
  wire al_60ceba51;
  wire al_763891b1;
  wire al_66ecf32f;
  wire al_cae9c79a;
  wire al_7fc110d7;
  wire al_26eaf94a;
  wire al_53f15a3f;
  wire al_ae71aa12;
  wire al_3f0ffcfa;
  wire al_d42a4c18;
  wire al_cf20ff1a;
  wire al_9ece8f02;
  wire al_8c6e2d36;
  wire al_3f77cd67;
  wire al_a8d42a04;
  wire al_388a24e;
  wire al_faa9857b;
  wire al_682de89f;
  wire al_f8ee3a1f;
  wire al_3d1ba91a;
  wire al_bdf8d79f;
  wire al_266f6c4c;
  wire al_f79b31c1;
  wire al_73642f31;
  wire al_7b4de920;
  wire al_b5c79ef6;
  wire al_87c0c365;
  wire al_9ba351db;
  wire al_eaafd789;
  wire al_100aadd6;
  wire al_38320d7c;
  wire al_1440c0b1;
  wire al_f6cc79fd;
  wire al_9ce6a803;
  wire al_4bdde34;
  wire al_6becface;
  wire al_136addab;
  wire al_c2479eab;
  wire al_c9c0fa32;
  wire al_c2428aac;
  wire al_8e6107a7;
  wire al_32c6ecc7;
  wire al_15bf91ee;
  wire al_d73f3ba1;
  wire al_af4842d7;
  wire al_336bd542;
  wire al_72f63008;
  wire al_5563a8fd;
  wire al_a51573d2;
  wire al_adae5a89;
  wire al_846b6533;
  wire al_9a1b441a;
  wire al_77e56b3a;
  wire al_807f5a12;
  wire al_7694b99f;
  wire al_3deafd60;
  wire al_67f58f23;
  wire al_c8a3ac58;
  wire al_46a6aa32;
  wire al_4ab17dc7;
  wire al_f718b05a;
  wire al_53f06a44;
  wire al_376757cc;
  wire al_83146215;
  wire al_c710cf1a;
  wire al_3d294c28;
  wire al_a5c6fbcc;
  wire al_cf358e1e;
  wire al_9aa134ca;
  wire al_e5bd99ae;
  wire al_e11118e;
  wire al_165ae4d7;
  wire al_8e1ef4c5;
  wire al_31ffb8d1;
  wire al_d0093be6;
  wire al_29396e02;
  wire al_e1b52e50;
  wire al_b05da9fd;
  wire al_160ccdf;
  wire al_a50584b2;
  wire al_c1b27879;
  wire al_803bd5d9;
  wire al_3daf6177;
  wire al_aa4375dc;
  wire al_f6a2d163;
  wire al_cd3c4af6;
  wire al_5ed94f60;
  wire al_db1fbb11;
  wire al_55ac2d11;
  wire al_d1cfb12d;
  wire al_f396fdd4;
  wire al_5a579dd;
  wire al_3e1dba29;
  wire al_5c82d563;
  wire al_a2faab7b;
  wire al_6f12ed1d;
  wire al_ef80f5cf;
  wire al_9b760ae7;
  wire al_290f1a7e;
  wire al_14c1cb65;
  wire al_32e957a5;
  wire al_b241735d;
  wire al_3fc75a33;
  wire al_e5994b5e;
  wire al_d8c8c74d;
  wire al_36c5508;
  wire al_5dda436f;
  wire al_c6a375ec;
  wire al_71ed2e0a;
  wire al_a78f40cd;
  wire al_78612548;
  wire al_64320b18;
  wire al_2162c82e;
  wire al_2c24255b;
  wire al_4ce1f25a;
  wire al_46d73024;
  wire al_b02bbd88;
  wire al_57b095a8;
  wire al_290af98f;
  wire al_7b30ef6a;
  wire al_870286f7;
  wire al_96ecb37f;
  wire al_482b5978;
  wire al_adc2de29;
  wire al_a2667927;
  wire al_efdbdafe;
  wire al_a8e6ffb8;
  wire al_35f24fff;
  wire al_ac79ddb;
  wire al_9e425de4;
  wire al_ebd2d7;
  wire al_857e17ab;
  wire al_7521303d;
  wire al_37168961;
  wire al_b48e2d4e;
  wire al_efc518d8;
  wire al_6b8a9b19;
  wire al_67b72f88;
  wire al_5ce38362;
  wire al_e0dc1ae0;
  wire al_762c3367;
  wire al_dcbb090f;
  wire al_153acd6e;
  wire al_94871a17;
  wire al_aa32962e;
  wire al_b96742e9;
  wire al_6f78b0c1;
  wire al_aaba7825;
  wire al_63eeda3d;
  wire al_76e16a6c;
  wire al_3fe47357;
  wire al_250851df;
  wire al_f5fd4d02;
  wire al_2d5ca5c8;
  wire al_765cb78c;
  wire al_618f3df7;
  wire al_9953d0c8;
  wire al_da48a386;
  wire al_3bac4202;
  wire al_27722f64;
  wire al_8c59fe48;
  wire al_bfd01551;
  wire al_fb3b1f47;
  wire al_fb660f65;
  wire al_c0e7d6fc;
  wire al_a381b363;
  wire al_84db8eae;
  wire al_27b5418b;
  wire al_de2d167c;
  wire al_da5e606a;
  wire al_f5fb13b0;
  wire al_f65615d7;
  wire al_fe5b64db;
  wire al_f3e72725;
  wire al_cd9f7a57;
  wire al_1717406d;
  wire al_74608a10;
  wire al_34e054a0;
  wire al_a3d91059;
  wire al_862844a1;
  wire al_62aa372c;
  wire al_6ed289d3;
  wire al_58e1cc88;
  wire al_e9ae3746;
  wire al_4a2b9f40;
  wire al_7c0f8e52;
  wire al_24faf4d6;
  wire al_5c9e751b;
  wire al_26e8cb8e;
  wire al_abe786cc;
  wire al_bd8e6c56;
  wire al_b1649623;
  wire al_4024362;
  wire al_496839d3;
  wire al_49948f6;
  wire al_783fafdc;
  wire al_a3ff8a2f;
  wire al_7f4e8532;
  wire al_12ae2ff1;
  wire al_f2f998df;
  wire al_f07e3782;
  wire al_6d77788f;
  wire al_b4f442b4;
  wire al_4c288bd1;
  wire al_232d54d1;
  wire al_465185e7;
  wire al_11d61e7f;
  wire al_ec82248c;
  wire al_130ad14e;
  wire al_e9c121e6;
  wire al_32e05e5d;
  wire al_d7d3035f;
  wire al_571ce91a;
  wire al_75707d25;
  wire al_abc33f01;
  wire al_8fda147c;
  wire al_c67dfcb5;
  wire al_ac325ba1;
  wire al_ebd48591;
  wire al_7b86230a;
  wire al_c98ce1a9;
  wire al_24ea5277;
  wire al_c560f884;
  wire al_8f7895f1;
  wire al_c198e7cb;
  wire al_bd399f0f;
  wire al_76c6b29d;
  wire al_cc7e8768;
  wire al_637261f7;
  wire al_aca9177e;
  wire al_f5473a34;
  wire al_69d9a189;
  wire al_be4e813d;
  wire al_c9ac0c17;
  wire al_cc5f5ce9;
  wire al_d0f70766;
  wire al_223a077f;
  wire al_db3a7a8b;
  wire al_297252e3;
  wire al_f44488cf;
  wire al_9e004fa1;
  wire al_5a460c8d;
  wire al_e7ad9386;
  wire al_f5f522a1;
  wire al_ab57e6bf;
  wire al_4cbbfdff;
  wire al_6300fa05;
  wire al_842395e3;
  wire al_69351137;
  wire al_514ce749;
  wire al_b04a4f00;
  wire al_5530c5c4;
  wire al_70e872b4;
  wire al_631f19c6;
  wire al_56607029;
  wire al_581760eb;
  wire al_b6529d32;
  wire al_53a5d1d8;
  wire al_263a3554;
  wire al_ccdce37d;
  wire al_ca35642e;
  wire al_5f4286cf;
  wire al_dcfb58ce;
  wire al_4276a847;
  wire al_a9c2861c;
  wire al_9daabc69;
  wire al_74d19130;
  wire al_a6104abc;
  wire al_271d4011;
  wire al_bd7f0fdb;
  wire al_1bd7127;
  wire al_4c1d19df;
  wire al_b42a6639;
  wire al_58a4ea01;
  wire al_c4d87e5a;
  wire al_56237b7;
  wire al_bf03de15;
  wire al_af6ff858;
  wire al_d50b6ef8;
  wire al_5f463be1;
  wire al_a927014c;
  wire al_acd7ad28;
  wire al_859e5564;
  wire al_772d3492;
  wire al_8a20aaa;
  wire al_b4bb4546;
  wire al_d2a71eb2;
  wire al_a2fcb15d;
  wire al_4d4393c7;
  wire al_d0651bd8;
  wire al_b77a14d7;
  wire al_8744257b;
  wire al_ded15eae;
  wire al_137e8f12;
  wire al_2408cdae;
  wire al_a63c88b4;
  wire al_83be6442;
  wire al_b0d20bea;
  wire al_98c88117;
  wire al_4a2c328a;
  wire al_ec1c3fd8;
  wire al_8c91da92;
  wire al_7f22fda0;
  wire al_8af9f67c;
  wire al_a808afa8;
  wire al_8a909a7e;
  wire al_7a2b8846;
  wire al_999473bf;
  wire al_3dc2993c;
  wire al_8e9644e7;
  wire al_54a9598a;
  wire al_85f33b95;
  wire al_c03c1e89;
  wire al_df93f3b6;
  wire al_bc71b143;
  wire al_c6d8833c;
  wire al_abb85d9;
  wire al_4503fb38;
  wire al_8298897d;
  wire al_56a26cfa;
  wire al_58887de;
  wire al_9073553b;
  wire al_d8b60780;
  wire al_4e2b6f95;
  wire al_513305d5;
  wire al_d7f7aaa1;
  wire al_c2044b3b;
  wire al_dbd06164;
  wire al_34ca3fbe;
  wire al_4f0b110;
  wire al_ac502f3b;
  wire al_b5cc7793;
  wire al_503c8f93;
  wire al_a81bacbe;
  wire al_72c24a7e;
  wire al_d67debd3;
  wire al_809052dd;
  wire al_6be58e65;
  wire al_95fe37a9;
  wire al_c8d005d;
  wire al_aacf80e2;
  wire al_68eb24f8;
  wire al_a07f4463;
  wire al_78627e02;
  wire al_bc4e38bd;
  wire al_96662c62;
  wire al_939c27b7;
  wire al_d9d7cf90;
  wire al_13db00fa;
  wire al_5bd0f2bc;
  wire al_484c4f9e;
  wire al_feb6df53;
  wire al_a3910e3c;
  wire al_3aba2254;
  wire al_51c4207;
  wire al_1855fcf8;
  wire al_855200e6;
  wire al_182d4638;
  wire al_63cbf333;
  wire al_63efbaa0;
  wire al_6e1ce9f;
  wire al_ae77f168;
  wire al_8213bac0;
  wire al_2b4ea789;
  wire al_9e8adc84;
  wire al_abdb8956;
  wire al_20628f76;

  assign gmii_tx_en = al_d32c67d0;
  assign gmii_tx_er = al_31529785;
  assign gmii_txd[7] = al_42702950[7];
  assign gmii_txd[6] = al_42702950[6];
  assign gmii_txd[5] = al_42702950[5];
  assign gmii_txd[4] = al_42702950[4];
  assign gmii_txd[3] = al_42702950[3];
  assign gmii_txd[2] = al_42702950[2];
  assign gmii_txd[1] = al_42702950[1];
  assign gmii_txd[0] = al_42702950[0];
  assign s_axi_bresp[1] = 1'b0;
  assign s_axi_bresp[0] = 1'b0;
  assign s_axi_rresp[1] = 1'b0;
  assign s_axi_rresp[0] = 1'b0;
  assign s_axi_wready = s_axi_awready;
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~A*~(D*C*~B)))"),
    .INIT(32'h0000baaa))
    al_2dca3acb (
    .a(tx_status_vector[3]),
    .b(al_67a4bdfd[0]),
    .c(al_67a4bdfd[1]),
    .d(al_67a4bdfd[4]),
    .e(tx_status_vld),
    .o(al_c9465832));
  AL_DFF_X al_acc6c02b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c9465832),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[3]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_17bd13d2 (
    .a(al_aeb75558[2]),
    .b(al_aeb75558[3]),
    .c(al_aeb75558[4]),
    .d(al_aeb75558[5]),
    .e(al_aeb75558[6]),
    .f(al_aeb75558[7]),
    .o(al_e18e0a15));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000010000))
    al_498c54a1 (
    .a(al_f6e00c9[4]),
    .b(al_f6e00c9[5]),
    .c(al_f6e00c9[6]),
    .d(al_f6e00c9[7]),
    .e(al_aeb75558[0]),
    .f(al_aeb75558[1]),
    .o(al_2de0dbf6));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_b9753c18 (
    .a(al_e18e0a15),
    .b(al_2de0dbf6),
    .c(al_f6e00c9[0]),
    .d(al_f6e00c9[1]),
    .e(al_f6e00c9[2]),
    .f(al_f6e00c9[3]),
    .o(al_c2be7784));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    al_4519b681 (
    .a(al_47e69606[0]),
    .b(al_47e69606[1]),
    .c(al_47e69606[2]),
    .d(al_47e69606[3]),
    .e(al_47e69606[4]),
    .o(al_a523c2cb));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~C*~(B*~A)))"),
    .INIT(32'h000000f4))
    al_a80b3a74 (
    .a(al_c2be7784),
    .b(al_a523c2cb),
    .c(al_4dabd984),
    .d(al_a37dea2d),
    .e(al_c99d4c23),
    .o(al_430719be));
  AL_DFF_X al_f1508bfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_430719be),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_4dabd984));
  AL_MAP_LUT6 #(
    .EQN("(A*~((E*~D*~C*B))*~(F)+A*(E*~D*~C*B)*~(F)+~(A)*~((E*~D*~C*B))*F)"),
    .INIT(64'h55515555aaaaaaaa))
    al_98f63a4d (
    .a(al_47e69606[0]),
    .b(al_47e69606[1]),
    .c(al_47e69606[2]),
    .d(al_47e69606[3]),
    .e(al_47e69606[4]),
    .f(al_c2520419),
    .o(al_a6a28e17[0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_43b9e7a9 (
    .a(al_a6a28e17[0]),
    .b(al_a37dea2d),
    .c(al_c99d4c23),
    .o(al_2b21b090[0]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~C*(B@(D*A)))"),
    .INIT(32'h0000060c))
    al_2ebda6d0 (
    .a(al_47e69606[0]),
    .b(al_47e69606[1]),
    .c(al_a37dea2d),
    .d(al_c2520419),
    .e(al_c99d4c23),
    .o(al_2b21b090[1]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~D*(C@(E*B*A)))"),
    .INIT(64'h00000000007800f0))
    al_b9ea9231 (
    .a(al_47e69606[0]),
    .b(al_47e69606[1]),
    .c(al_47e69606[2]),
    .d(al_a37dea2d),
    .e(al_c2520419),
    .f(al_c99d4c23),
    .o(al_2b21b090[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*C*B*A))"),
    .INIT(32'h7f80ff00))
    al_60cf3b13 (
    .a(al_47e69606[0]),
    .b(al_47e69606[1]),
    .c(al_47e69606[2]),
    .d(al_47e69606[3]),
    .e(al_c2520419),
    .o(al_a6a28e17[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_22b273f0 (
    .a(al_a6a28e17[3]),
    .b(al_a37dea2d),
    .c(al_c99d4c23),
    .o(al_2b21b090[3]));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*D*C*B*A))"),
    .INIT(64'h7fff8000ffff0000))
    al_58b009e (
    .a(al_47e69606[0]),
    .b(al_47e69606[1]),
    .c(al_47e69606[2]),
    .d(al_47e69606[3]),
    .e(al_47e69606[4]),
    .f(al_c2520419),
    .o(al_a6a28e17[4]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_e70346e5 (
    .a(al_a6a28e17[4]),
    .b(al_a37dea2d),
    .c(al_c99d4c23),
    .o(al_2b21b090[4]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~C*~(B*A)))"),
    .INIT(32'h000000f8))
    al_d29a65f9 (
    .a(al_c2be7784),
    .b(al_a523c2cb),
    .c(al_b2b271cb),
    .d(al_a37dea2d),
    .e(al_c99d4c23),
    .o(al_4d9c2a7a));
  AL_DFF_X al_b7d0217d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4d9c2a7a),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_b2b271cb));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_d63c89f4 (
    .a(al_5a6020b4),
    .b(al_e1f88382[0]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[0]),
    .o(al_e6e0b636[0]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_cf911c70 (
    .a(al_82120dcc),
    .b(al_e1f88382[10]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[2]),
    .o(al_e6e0b636[10]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_2333dd2e (
    .a(al_82120dcc),
    .b(al_e1f88382[11]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[3]),
    .o(al_e6e0b636[11]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_ca87d2aa (
    .a(al_82120dcc),
    .b(al_e1f88382[12]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[4]),
    .o(al_e6e0b636[12]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_510fd775 (
    .a(al_82120dcc),
    .b(al_e1f88382[13]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[5]),
    .o(al_e6e0b636[13]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_b962fad7 (
    .a(al_82120dcc),
    .b(al_e1f88382[14]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[6]),
    .o(al_e6e0b636[14]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    al_3e128455 (
    .a(al_47e69606[0]),
    .b(al_47e69606[1]),
    .c(al_47e69606[2]),
    .d(al_47e69606[3]),
    .e(al_47e69606[4]),
    .o(al_82120dcc));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_458d36ee (
    .a(al_82120dcc),
    .b(al_e1f88382[15]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[7]),
    .o(al_e6e0b636[15]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_2893dfbf (
    .a(al_5a6020b4),
    .b(al_e1f88382[1]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[1]),
    .o(al_e6e0b636[1]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_793860ae (
    .a(al_5a6020b4),
    .b(al_e1f88382[2]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[2]),
    .o(al_e6e0b636[2]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_cda8bdd7 (
    .a(al_5a6020b4),
    .b(al_e1f88382[3]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[3]),
    .o(al_e6e0b636[3]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_fc7cc981 (
    .a(al_5a6020b4),
    .b(al_e1f88382[4]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[4]),
    .o(al_e6e0b636[4]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_69cbe49f (
    .a(al_5a6020b4),
    .b(al_e1f88382[5]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[5]),
    .o(al_e6e0b636[5]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_c46740ac (
    .a(al_5a6020b4),
    .b(al_e1f88382[6]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[6]),
    .o(al_e6e0b636[6]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_f8f10ac7 (
    .a(al_47e69606[0]),
    .b(al_47e69606[1]),
    .c(al_47e69606[2]),
    .d(al_47e69606[3]),
    .e(al_47e69606[4]),
    .o(al_5a6020b4));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_67fe4ec9 (
    .a(al_5a6020b4),
    .b(al_e1f88382[7]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[7]),
    .o(al_e6e0b636[7]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_1452da83 (
    .a(al_82120dcc),
    .b(al_e1f88382[8]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[0]),
    .o(al_e6e0b636[8]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(B*~(E)*~(A)+B*E*~(A)+~(B)*E*A+B*E*A))"),
    .INIT(32'h000e0004))
    al_9cebad15 (
    .a(al_82120dcc),
    .b(al_e1f88382[9]),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_aeb75558[1]),
    .o(al_e6e0b636[9]));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*D*C*~B*A)"),
    .INIT(64'h0000000020000000))
    al_c6ea618f (
    .a(rx_clk_en),
    .b(al_47e69606[0]),
    .c(al_47e69606[1]),
    .d(al_47e69606[2]),
    .e(al_47e69606[3]),
    .f(al_47e69606[4]),
    .o(al_a6ff135b));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_f5de3a2b (
    .a(al_a6ff135b),
    .b(al_a37dea2d),
    .c(al_c99d4c23),
    .o(al_aaead9c7));
  AL_DFF_X al_61486ff5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2b21b090[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_47e69606[0]));
  AL_DFF_X al_9c157454 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2b21b090[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_47e69606[1]));
  AL_DFF_X al_912d724c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2b21b090[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_47e69606[2]));
  AL_DFF_X al_c073d488 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2b21b090[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_47e69606[3]));
  AL_DFF_X al_6b613f07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2b21b090[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_47e69606[4]));
  AL_DFF_X al_e95068a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[0]),
    .en(al_aaead9c7),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f6e00c9[0]));
  AL_DFF_X al_70b53be7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[1]),
    .en(al_aaead9c7),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f6e00c9[1]));
  AL_DFF_X al_ac801176 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[2]),
    .en(al_aaead9c7),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f6e00c9[2]));
  AL_DFF_X al_fbd81f4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[3]),
    .en(al_aaead9c7),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f6e00c9[3]));
  AL_DFF_X al_afe3b421 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[4]),
    .en(al_aaead9c7),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f6e00c9[4]));
  AL_DFF_X al_65eb47bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[5]),
    .en(al_aaead9c7),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f6e00c9[5]));
  AL_DFF_X al_99b32eb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[6]),
    .en(al_aaead9c7),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f6e00c9[6]));
  AL_DFF_X al_2cd98aef (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[7]),
    .en(al_aaead9c7),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f6e00c9[7]));
  AL_DFF_X al_718a4ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[8]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[8]));
  AL_DFF_X al_76de083d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[9]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[9]));
  AL_DFF_X al_9eb34218 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[10]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[10]));
  AL_DFF_X al_61f97cbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[11]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[11]));
  AL_DFF_X al_dae5b7c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[12]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[12]));
  AL_DFF_X al_632bc37a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[13]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[13]));
  AL_DFF_X al_7bd43bf8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[14]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[14]));
  AL_DFF_X al_f7d071ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[15]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[15]));
  AL_DFF_X al_e2a63491 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[0]));
  AL_DFF_X al_94498507 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[1]));
  AL_DFF_X al_ddd84bbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[2]));
  AL_DFF_X al_43d59b2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[3]));
  AL_DFF_X al_21b4f197 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[4]));
  AL_DFF_X al_d93fe8ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[5]));
  AL_DFF_X al_c5ba0c59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[6]));
  AL_DFF_X al_76c5f02c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e6e0b636[7]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1f88382[7]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(E*D*~B*A))"),
    .INIT(32'hf2f0f0f0))
    al_a3919ab0 (
    .a(al_6bdd801e),
    .b(al_4dabd984),
    .c(al_a37dea2d),
    .d(al_c99d4c23),
    .e(al_b2deb19c),
    .o(al_5b289734));
  AL_DFF_X al_7afd9215 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5b289734),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_error_frame));
  AL_DFF_X al_8f1cd930 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c2520419),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_data_vld));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d0fcef1d (
    .a(al_e495ee45),
    .b(al_a76fca28),
    .o(al_f164e0a));
  AL_DFF_X al_7cfab1ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f164e0a),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_6bdd801e));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~B*A))"),
    .INIT(16'hd0f0))
    al_91262812 (
    .a(al_6bdd801e),
    .b(al_4dabd984),
    .c(al_c99d4c23),
    .d(al_b2deb19c),
    .o(al_74354c6e));
  AL_DFF_X al_f3b1bc0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_74354c6e),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_correct_frame));
  AL_DFF_X al_a5cba89b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c99d4c23),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_93abd71));
  AL_DFF_X al_22728197 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_93abd71),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_3a74e04b));
  AL_DFF_X al_bcb3ad8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_3a74e04b),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_33e46ce3));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_29a07068 (
    .a(al_93abd71),
    .b(al_3a74e04b),
    .c(al_33e46ce3),
    .o(al_6b96fb99));
  AL_DFF_X al_6995a34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6b96fb99),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_47f8fdc1));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_e4db5359 (
    .a(rx_clk_en),
    .b(al_c99d4c23),
    .o(al_18e5b9af));
  AL_DFF_X al_3788d16c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_51616140),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f55c93aa));
  AL_DFF_X al_169032b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[8]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[8]));
  AL_DFF_X al_34e6980a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[9]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[9]));
  AL_DFF_X al_43986354 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[10]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[10]));
  AL_DFF_X al_fca65d9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[11]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[11]));
  AL_DFF_X al_b96db99e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[12]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[12]));
  AL_DFF_X al_e11f3a23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[13]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[13]));
  AL_DFF_X al_d6ce665 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[14]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[14]));
  AL_DFF_X al_d68c4330 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[15]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[15]));
  AL_DFF_X al_d1ba941d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[0]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[0]));
  AL_DFF_X al_d1ca4c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[1]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[1]));
  AL_DFF_X al_d3ff55ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[2]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[2]));
  AL_DFF_X al_1726dd92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[3]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[3]));
  AL_DFF_X al_8f809105 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[4]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[4]));
  AL_DFF_X al_69f619aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[5]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[5]));
  AL_DFF_X al_95003808 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[6]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[6]));
  AL_DFF_X al_f7cde603 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1f88382[7]),
    .en(al_18e5b9af),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7d74a9c[7]));
  AL_DFF_X al_4aeb4350 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1440c0b1),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_b65ba3d5));
  AL_DFF_X al_54a493dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1bba34ee),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9eb158b7));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_d82fd82b (
    .a(tx_data_en),
    .b(al_9eb158b7),
    .o(tx_rdy));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_ce7f9302 (
    .a(al_9953d0c8),
    .b(al_2a1554ab[0]),
    .c(al_2a1554ab[1]),
    .d(al_2a1554ab[2]),
    .o(al_1440c0b1));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~B*~(~D*C*A)))"),
    .INIT(32'h0000ccec))
    al_1a6bf9cd (
    .a(al_1440c0b1),
    .b(tx_rdy),
    .c(tx_clk_en),
    .d(al_7dd23876),
    .e(al_2dbca608),
    .o(al_1bba34ee));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~((~E*~D*~C))*~(F)+(~B*~A)*~((~E*~D*~C))*~(F)+~((~B*~A))*(~E*~D*~C)*~(F)+~((~B*~A))*(~E*~D*~C)*F+(~B*~A)*(~E*~D*~C)*F)"),
    .INIT(64'h0000000ffffffffe))
    al_44fccf82 (
    .a(al_d1c7d2fd),
    .b(al_67a4bdfd[0]),
    .c(al_67a4bdfd[1]),
    .d(al_67a4bdfd[2]),
    .e(al_67a4bdfd[3]),
    .f(al_67a4bdfd[4]),
    .o(al_d7389040));
  AL_DFF_X al_c27142e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d7389040),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1421d0c8));
  AL_DFF_X al_3abc778e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data_en),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_ac2b4841));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_c9f0ebeb (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_c5235ca5[16]),
    .d(al_c5235ca5[24]),
    .e(al_c5235ca5[32]),
    .f(al_c5235ca5[40]),
    .o(al_1da67580));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fd264819 (
    .a(al_67a4bdfd[0]),
    .b(al_c5235ca5[0]),
    .c(al_c5235ca5[8]),
    .o(al_bf066204));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F)"),
    .INIT(64'h0fffaaaa330ffff0))
    al_4c957bc5 (
    .a(al_1da67580),
    .b(al_bf066204),
    .c(al_67a4bdfd[0]),
    .d(al_67a4bdfd[1]),
    .e(al_67a4bdfd[2]),
    .f(al_67a4bdfd[3]),
    .o(al_889a47a2));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hcd458901))
    al_1e54cd58 (
    .a(al_889a47a2),
    .b(al_e2a1fab3),
    .c(al_67a4bdfd[4]),
    .d(al_522cbac[0]),
    .e(al_522cbac[8]),
    .o(al_de1356f0[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_897c3fd9 (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_c5235ca5[17]),
    .d(al_c5235ca5[25]),
    .e(al_c5235ca5[33]),
    .f(al_c5235ca5[41]),
    .o(al_65719225));
  AL_MAP_LUT5 #(
    .EQN("(B*(~(A)*~(C)*~(D)*~(E)+~(A)*~(C)*D*~(E)+~(A)*C*D*~(E)+~(A)*~(C)*~(D)*E+A*C*~(D)*E+~(A)*~(C)*D*E+~(A)*C*D*E+A*C*D*E))"),
    .INIT(32'hc4844404))
    al_117e563a (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_67a4bdfd[2]),
    .d(al_c5235ca5[1]),
    .e(al_c5235ca5[9]),
    .o(al_de41ced));
  AL_MAP_LUT5 #(
    .EQN("(~E*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .INIT(32'h000005cc))
    al_4cbc748d (
    .a(al_65719225),
    .b(al_de41ced),
    .c(al_67a4bdfd[2]),
    .d(al_67a4bdfd[3]),
    .e(al_67a4bdfd[4]),
    .o(al_5d511a0d));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(B*(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)))"),
    .INIT(32'heeaeeaaa))
    al_69c981c2 (
    .a(al_5d511a0d),
    .b(al_e2a1fab3),
    .c(al_67a4bdfd[0]),
    .d(al_522cbac[1]),
    .e(al_522cbac[9]),
    .o(al_de1356f0[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_e07ea270 (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_c5235ca5[18]),
    .d(al_c5235ca5[26]),
    .e(al_c5235ca5[34]),
    .f(al_c5235ca5[42]),
    .o(al_1a69e04c));
  AL_MAP_LUT6 #(
    .EQN("(~((E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D)*B)*~(C*~A))"),
    .INIT(64'h232323afaf23afaf))
    al_f062e05d (
    .a(al_1a69e04c),
    .b(al_90044ea4),
    .c(al_4b956df0),
    .d(al_67a4bdfd[0]),
    .e(al_c5235ca5[2]),
    .f(al_c5235ca5[10]),
    .o(al_4940717b));
  AL_MAP_LUT6 #(
    .EQN("~(~((F*~(E)*~(C)+F*E*~(C)+~(F)*E*C+F*E*C)*B)*~(~D*~A))"),
    .INIT(64'hccdd0c5dc0d50055))
    al_e86c2cc3 (
    .a(al_4940717b),
    .b(al_e2a1fab3),
    .c(al_67a4bdfd[0]),
    .d(al_67a4bdfd[4]),
    .e(al_522cbac[2]),
    .f(al_522cbac[10]),
    .o(al_de1356f0[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_68d4f9a6 (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_c5235ca5[19]),
    .d(al_c5235ca5[27]),
    .e(al_c5235ca5[35]),
    .f(al_c5235ca5[43]),
    .o(al_abceb3af));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_88332102 (
    .a(al_67a4bdfd[0]),
    .b(al_c5235ca5[3]),
    .c(al_c5235ca5[11]),
    .o(al_76834e7a));
  AL_MAP_LUT6 #(
    .EQN("(~F*(~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E))"),
    .INIT(64'h000000000f55c000))
    al_3df769f4 (
    .a(al_abceb3af),
    .b(al_76834e7a),
    .c(al_67a4bdfd[1]),
    .d(al_67a4bdfd[2]),
    .e(al_67a4bdfd[3]),
    .f(al_67a4bdfd[4]),
    .o(al_d9c2bbe5));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(B*(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)))"),
    .INIT(32'heeaeeaaa))
    al_ef5876a4 (
    .a(al_d9c2bbe5),
    .b(al_e2a1fab3),
    .c(al_67a4bdfd[0]),
    .d(al_522cbac[3]),
    .e(al_522cbac[11]),
    .o(al_de1356f0[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_40ae7153 (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_c5235ca5[20]),
    .d(al_c5235ca5[28]),
    .e(al_c5235ca5[36]),
    .f(al_c5235ca5[44]),
    .o(al_b93d302f));
  AL_MAP_LUT6 #(
    .EQN("(~((E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D)*B)*~(C*~A))"),
    .INIT(64'h232323afaf23afaf))
    al_677952b8 (
    .a(al_b93d302f),
    .b(al_90044ea4),
    .c(al_4b956df0),
    .d(al_67a4bdfd[0]),
    .e(al_c5235ca5[4]),
    .f(al_c5235ca5[12]),
    .o(al_fd543856));
  AL_MAP_LUT6 #(
    .EQN("~(~((F*~(E)*~(C)+F*E*~(C)+~(F)*E*C+F*E*C)*B)*~(~D*~A))"),
    .INIT(64'hccdd0c5dc0d50055))
    al_72405bd8 (
    .a(al_fd543856),
    .b(al_e2a1fab3),
    .c(al_67a4bdfd[0]),
    .d(al_67a4bdfd[4]),
    .e(al_522cbac[4]),
    .f(al_522cbac[12]),
    .o(al_de1356f0[4]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_7f6063b9 (
    .a(al_67a4bdfd[1]),
    .b(al_67a4bdfd[2]),
    .c(al_67a4bdfd[3]),
    .o(al_90044ea4));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_9796e9a0 (
    .a(al_67a4bdfd[2]),
    .b(al_67a4bdfd[3]),
    .o(al_4b956df0));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_b42c8344 (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_c5235ca5[21]),
    .d(al_c5235ca5[29]),
    .e(al_c5235ca5[37]),
    .f(al_c5235ca5[45]),
    .o(al_a88739b8));
  AL_MAP_LUT6 #(
    .EQN("(~((E*~(F)*~(D)+E*F*~(D)+~(E)*F*D+E*F*D)*B)*~(C*~A))"),
    .INIT(64'h232323afaf23afaf))
    al_61ed3f99 (
    .a(al_a88739b8),
    .b(al_90044ea4),
    .c(al_4b956df0),
    .d(al_67a4bdfd[0]),
    .e(al_c5235ca5[5]),
    .f(al_c5235ca5[13]),
    .o(al_eeb871e3));
  AL_MAP_LUT6 #(
    .EQN("~(~((F*~(E)*~(C)+F*E*~(C)+~(F)*E*C+F*E*C)*B)*~(~D*~A))"),
    .INIT(64'hccdd0c5dc0d50055))
    al_f15d8ea1 (
    .a(al_eeb871e3),
    .b(al_e2a1fab3),
    .c(al_67a4bdfd[0]),
    .d(al_67a4bdfd[4]),
    .e(al_522cbac[5]),
    .f(al_522cbac[13]),
    .o(al_de1356f0[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_40bd7165 (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_c5235ca5[22]),
    .d(al_c5235ca5[30]),
    .e(al_c5235ca5[38]),
    .f(al_c5235ca5[46]),
    .o(al_c192e229));
  AL_MAP_LUT5 #(
    .EQN("(B*(~(A)*~(C)*~(D)*~(E)+~(A)*~(C)*D*~(E)+~(A)*C*D*~(E)+~(A)*~(C)*~(D)*E+A*C*~(D)*E+~(A)*~(C)*D*E+~(A)*C*D*E+A*C*D*E))"),
    .INIT(32'hc4844404))
    al_78e811ca (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_67a4bdfd[2]),
    .d(al_c5235ca5[6]),
    .e(al_c5235ca5[14]),
    .o(al_84a2caa3));
  AL_MAP_LUT5 #(
    .EQN("(~E*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .INIT(32'h000005cc))
    al_9290529d (
    .a(al_c192e229),
    .b(al_84a2caa3),
    .c(al_67a4bdfd[2]),
    .d(al_67a4bdfd[3]),
    .e(al_67a4bdfd[4]),
    .o(al_5ecede8f));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(B*(E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)))"),
    .INIT(32'heeaeeaaa))
    al_349b0d14 (
    .a(al_5ecede8f),
    .b(al_e2a1fab3),
    .c(al_67a4bdfd[0]),
    .d(al_522cbac[6]),
    .e(al_522cbac[14]),
    .o(al_de1356f0[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    al_d629f0aa (
    .a(al_67a4bdfd[1]),
    .b(al_67a4bdfd[2]),
    .c(al_67a4bdfd[3]),
    .d(al_67a4bdfd[4]),
    .o(al_e2a1fab3));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_cf25c77f (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_c5235ca5[23]),
    .d(al_c5235ca5[31]),
    .e(al_c5235ca5[39]),
    .f(al_c5235ca5[47]),
    .o(al_511fc342));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_334d6027 (
    .a(al_67a4bdfd[0]),
    .b(al_c5235ca5[7]),
    .c(al_c5235ca5[15]),
    .o(al_cba22e49));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff0aaaa33fff00f))
    al_1407bd27 (
    .a(al_511fc342),
    .b(al_cba22e49),
    .c(al_67a4bdfd[0]),
    .d(al_67a4bdfd[1]),
    .e(al_67a4bdfd[2]),
    .f(al_67a4bdfd[3]),
    .o(al_7f616b69));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hcd894501))
    al_24031bd3 (
    .a(al_7f616b69),
    .b(al_e2a1fab3),
    .c(al_67a4bdfd[4]),
    .d(al_522cbac[7]),
    .e(al_522cbac[15]),
    .o(al_de1356f0[7]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_4d46c71d (
    .a(al_69e62d6a),
    .b(al_f4206233),
    .c(al_67a4bdfd[0]),
    .o(al_cade1083[0]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ba0))
    al_f6061a2c (
    .a(al_69e62d6a),
    .b(al_f4206233),
    .c(al_67a4bdfd[0]),
    .d(al_67a4bdfd[1]),
    .o(al_cade1083[1]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*(D*C)*~(E)+A*B*(D*C)*~(E)+~(A)*~(B)*~((D*C))*E+A*~(B)*~((D*C))*E+A*B*~((D*C))*E+~(A)*~(B)*(D*C)*E)"),
    .INIT(32'h1bbba000))
    al_9a0164f (
    .a(al_69e62d6a),
    .b(al_f4206233),
    .c(al_67a4bdfd[0]),
    .d(al_67a4bdfd[1]),
    .e(al_67a4bdfd[2]),
    .o(al_cade1083[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*(E*D*C)*~(F)+A*B*(E*D*C)*~(F)+~(A)*~(B)*~((E*D*C))*F+A*~(B)*~((E*D*C))*F+A*B*~((E*D*C))*F+~(A)*~(B)*(E*D*C)*F)"),
    .INIT(64'h1bbbbbbba0000000))
    al_cec978fd (
    .a(al_69e62d6a),
    .b(al_f4206233),
    .c(al_67a4bdfd[0]),
    .d(al_67a4bdfd[1]),
    .e(al_67a4bdfd[2]),
    .f(al_67a4bdfd[3]),
    .o(al_cade1083[3]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    al_a376f56 (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_67a4bdfd[2]),
    .d(al_67a4bdfd[3]),
    .e(al_67a4bdfd[4]),
    .o(al_b306469e));
  AL_MAP_LUT5 #(
    .EQN("(D*C*~A*~(~E*~B))"),
    .INIT(32'h50004000))
    al_961f8e75 (
    .a(al_b306469e),
    .b(al_b65ba3d5),
    .c(al_7dd23876),
    .d(al_f4206233),
    .e(al_520772a3[2]),
    .o(al_69e62d6a));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_bb720146 (
    .a(al_67a4bdfd[0]),
    .b(al_67a4bdfd[1]),
    .c(al_67a4bdfd[2]),
    .d(al_67a4bdfd[3]),
    .o(al_82835dec));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h2f88))
    al_3f5ed0e5 (
    .a(al_69e62d6a),
    .b(al_82835dec),
    .c(al_f4206233),
    .d(al_67a4bdfd[4]),
    .o(al_cade1083[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    al_5edb8402 (
    .a(al_95c95cdd),
    .b(al_ac2b4841),
    .c(al_5e18973f),
    .o(al_fe501ed1));
  AL_DFF_X al_f283f293 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_fe501ed1),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_5e18973f));
  AL_DFF_X al_5c91ad71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_95c95cdd),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_d1c7d2fd));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*~B*A)"),
    .INIT(16'hdfff))
    al_98e0cbc2 (
    .a(al_73bb0740),
    .b(al_f79b31c1),
    .c(al_266f6c4c),
    .d(al_a381b363),
    .o(al_95c95cdd));
  AL_MAP_LUT5 #(
    .EQN("(B*~A*~(E*~D*~C))"),
    .INIT(32'h44404444))
    al_f5b1e014 (
    .a(al_f4206233),
    .b(al_520772a3[0]),
    .c(al_520772a3[1]),
    .d(al_520772a3[2]),
    .e(al_452dacc5),
    .o(al_a655b507));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~(A*~(C*B))))"),
    .INIT(32'h00002aff))
    al_a7df681a (
    .a(al_a655b507),
    .b(al_ac2b4841),
    .c(al_5e18973f),
    .d(al_7dd23876),
    .e(al_23e59594),
    .o(al_758baf6a));
  AL_MAP_LUT5 #(
    .EQN("~(A*~(~(~E*~D)*~(C*B)))"),
    .INIT(32'h7f7f7f55))
    al_159d6a53 (
    .a(al_758baf6a),
    .b(al_95c95cdd),
    .c(al_ac2b4841),
    .d(al_f4206233),
    .e(al_452dacc5),
    .o(al_b3b32038));
  AL_DFF_X al_90c58b8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b3b32038),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_7dd23876));
  AL_MAP_LUT6 #(
    .EQN("(~(F*E*~D)*~(~C*~(B*A)))"),
    .INIT(64'hf800f8f8f8f8f8f8))
    al_19ca88b4 (
    .a(pause_req),
    .b(al_c292362f),
    .c(al_f4206233),
    .d(al_67a4bdfd[0]),
    .e(al_67a4bdfd[1]),
    .f(al_67a4bdfd[4]),
    .o(al_82c4c889));
  AL_DFF_X al_f3bda375 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_82c4c889),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f4206233));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(A*~(E*D*~C)))"),
    .INIT(32'h13111111))
    al_4949cd9c (
    .a(al_ac2b4841),
    .b(al_7dd23876),
    .c(al_f79b31c1),
    .d(al_266f6c4c),
    .e(al_a381b363),
    .o(al_1c26630b));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~A*~(D*C*~B))"),
    .INIT(64'h0000455500000000))
    al_19e11757 (
    .a(al_1c26630b),
    .b(al_67a4bdfd[0]),
    .c(al_67a4bdfd[1]),
    .d(al_67a4bdfd[4]),
    .e(al_520772a3[1]),
    .f(al_520772a3[2]),
    .o(al_d78ef14f));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~A*~(~E*D*B)))"),
    .INIT(32'h0a0a0e0a))
    al_49d4ffb7 (
    .a(al_d78ef14f),
    .b(al_b65ba3d5),
    .c(al_520772a3[0]),
    .d(al_520772a3[1]),
    .e(al_520772a3[2]),
    .o(al_a51041a6));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~C*~B*A))"),
    .INIT(32'h00ff00fd))
    al_bc7ba151 (
    .a(al_ac2b4841),
    .b(al_5e18973f),
    .c(al_7dd23876),
    .d(al_f4206233),
    .e(al_23e59594),
    .o(al_5097d6f));
  AL_MAP_LUT5 #(
    .EQN("(~E*(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D))"),
    .INIT(32'h00000350))
    al_ed0a5056 (
    .a(al_5097d6f),
    .b(al_b65ba3d5),
    .c(al_520772a3[0]),
    .d(al_520772a3[1]),
    .e(al_520772a3[2]),
    .o(al_7fd108f9));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hf5f5f0c5))
    al_544214e (
    .a(al_d78ef14f),
    .b(al_5097d6f),
    .c(al_520772a3[0]),
    .d(al_520772a3[1]),
    .e(al_520772a3[2]),
    .o(al_6aba2287));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_6df2e56f (
    .a(tx_clk_en),
    .b(al_f4206233),
    .c(al_520772a3[0]),
    .o(al_eb74cd21));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_df86d552 (
    .a(pause_req),
    .b(tx_clk_en),
    .o(al_fb8448e4));
  AL_DFF_X al_f269f5db (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_de1356f0[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9c49a375[0]));
  AL_DFF_X al_b2192d43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_de1356f0[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9c49a375[1]));
  AL_DFF_X al_f7c66e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_de1356f0[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9c49a375[2]));
  AL_DFF_X al_ec7c0278 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_de1356f0[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9c49a375[3]));
  AL_DFF_X al_c3618feb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_de1356f0[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9c49a375[4]));
  AL_DFF_X al_26509d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_de1356f0[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9c49a375[5]));
  AL_DFF_X al_91bd3b43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_de1356f0[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9c49a375[6]));
  AL_DFF_X al_6ebda7d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_de1356f0[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9c49a375[7]));
  AL_DFF_X al_985f4024 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cade1083[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_67a4bdfd[0]));
  AL_DFF_X al_fb8d7299 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cade1083[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_67a4bdfd[1]));
  AL_DFF_X al_6b3da532 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cade1083[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_67a4bdfd[2]));
  AL_DFF_X al_b54ba2a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cade1083[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_67a4bdfd[3]));
  AL_DFF_X al_6ae16e7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cade1083[4]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_67a4bdfd[4]));
  AL_DFF_X al_a39ffadb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[8]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[8]));
  AL_DFF_X al_6a610256 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[9]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[9]));
  AL_DFF_X al_cff2e777 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[10]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[10]));
  AL_DFF_X al_a80f157d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[11]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[11]));
  AL_DFF_X al_ce576fb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[12]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[12]));
  AL_DFF_X al_5dab8417 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[13]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[13]));
  AL_DFF_X al_26a6ab71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[14]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[14]));
  AL_DFF_X al_418aa737 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[15]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[15]));
  AL_DFF_X al_d2d798bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[16]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[16]));
  AL_DFF_X al_7df8b19b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[17]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[17]));
  AL_DFF_X al_779065b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[0]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[0]));
  AL_DFF_X al_7ccb4a7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[18]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[18]));
  AL_DFF_X al_ca34cfee (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[19]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[19]));
  AL_DFF_X al_745cc8b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[20]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[20]));
  AL_DFF_X al_f59a09cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[21]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[21]));
  AL_DFF_X al_279bd9a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[22]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[22]));
  AL_DFF_X al_902f2b1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[23]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[23]));
  AL_DFF_X al_fb817561 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[24]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[24]));
  AL_DFF_X al_b35f1827 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[25]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[25]));
  AL_DFF_X al_303d7f52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[26]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[26]));
  AL_DFF_X al_77fab6f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[27]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[27]));
  AL_DFF_X al_5b30cf11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[1]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[1]));
  AL_DFF_X al_cae7e72d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[28]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[28]));
  AL_DFF_X al_360b020a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[29]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[29]));
  AL_DFF_X al_be27dbb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[30]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[30]));
  AL_DFF_X al_95b3477 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[31]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[31]));
  AL_DFF_X al_3329f864 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[0]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[32]));
  AL_DFF_X al_7f3b194f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[1]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[33]));
  AL_DFF_X al_712ca633 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[2]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[34]));
  AL_DFF_X al_c6e4fddd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[3]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[35]));
  AL_DFF_X al_1fd6bb4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[4]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[36]));
  AL_DFF_X al_65ffb5e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[5]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[37]));
  AL_DFF_X al_e0db744c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[2]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[2]));
  AL_DFF_X al_88afbb9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[6]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[38]));
  AL_DFF_X al_773264b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[7]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[39]));
  AL_DFF_X al_f60375a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[8]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[40]));
  AL_DFF_X al_e2e2567e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[9]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[41]));
  AL_DFF_X al_b78d95d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[10]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[42]));
  AL_DFF_X al_384e725c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[11]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[43]));
  AL_DFF_X al_dc4a9561 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[12]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[44]));
  AL_DFF_X al_812e18aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[13]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[45]));
  AL_DFF_X al_eb58ff25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[14]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[46]));
  AL_DFF_X al_9ec4458e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3c2ad2a[15]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[47]));
  AL_DFF_X al_8f4c728 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[3]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[3]));
  AL_DFF_X al_66b3b06f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[4]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[4]));
  AL_DFF_X al_b04de7c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[5]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[5]));
  AL_DFF_X al_4672fd3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[6]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[6]));
  AL_DFF_X al_9e4910b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_42381c95[7]),
    .en(al_eb74cd21),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5235ca5[7]));
  AL_DFF_X al_684c63b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[8]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[8]));
  AL_DFF_X al_737177b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[9]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[9]));
  AL_DFF_X al_98a9fc04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[10]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[10]));
  AL_DFF_X al_32aa3071 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[11]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[11]));
  AL_DFF_X al_2e19fca (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[12]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[12]));
  AL_DFF_X al_b3ef5359 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[13]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[13]));
  AL_DFF_X al_a16c025a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[14]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[14]));
  AL_DFF_X al_c5be39c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[15]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[15]));
  AL_DFF_X al_d6baea51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[0]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[0]));
  AL_DFF_X al_fc388eed (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[1]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[1]));
  AL_DFF_X al_2256c2fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[2]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[2]));
  AL_DFF_X al_2802e5ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[3]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[3]));
  AL_DFF_X al_d1e35682 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[4]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[4]));
  AL_DFF_X al_ca934a9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[5]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[5]));
  AL_DFF_X al_f04d606e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[6]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[6]));
  AL_DFF_X al_42a0352e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[7]),
    .en(al_fb8448e4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_522cbac[7]));
  AL_DFF_X al_2af1cb49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6aba2287),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_520772a3[0]));
  AL_DFF_X al_3c2b5424 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7fd108f9),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_520772a3[1]));
  AL_DFF_X al_e5b83089 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a51041a6),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_520772a3[2]));
  AL_DFF_X al_3021a46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5c82d563),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_collision));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_253e0474 (
    .a(al_715e8e22),
    .b(al_637ddda1),
    .o(al_5b37fe28));
  AL_DFF_X al_51c99fd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5b37fe28),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c292362f));
  AL_DFF_X al_416fd896 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_452dacc5),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9cae7666));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_87415e4e (
    .a(al_7d74a9c[10]),
    .b(al_7d74a9c[11]),
    .c(al_7d74a9c[12]),
    .d(al_7d74a9c[13]),
    .e(al_7d74a9c[14]),
    .f(al_7d74a9c[15]),
    .o(al_d811a788));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_70ac31c8 (
    .a(al_7d74a9c[4]),
    .b(al_7d74a9c[5]),
    .c(al_7d74a9c[6]),
    .d(al_7d74a9c[7]),
    .e(al_7d74a9c[8]),
    .f(al_7d74a9c[9]),
    .o(al_8e5a365f));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_f4ca99bb (
    .a(al_d811a788),
    .b(al_8e5a365f),
    .c(al_7d74a9c[0]),
    .d(al_7d74a9c[1]),
    .e(al_7d74a9c[2]),
    .f(al_7d74a9c[3]),
    .o(al_2c74b50c));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*C)*~(A)*~(B)+~(~D*C)*A*~(B)+~(~(~D*C))*A*B+~(~D*C)*A*B)"),
    .INIT(16'h4474))
    al_c4e345e9 (
    .a(al_2c74b50c),
    .b(al_c92c521a),
    .c(al_452dacc5),
    .d(al_23e59594),
    .o(al_495ac57d));
  AL_DFF_X al_3225b512 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_495ac57d),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_452dacc5));
  AL_DFF_X al_99497a5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6127633d),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f9514cde));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_1e3f7b43 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[0]),
    .d(al_64a46519[0]),
    .e(al_8a4cc919[0]),
    .o(al_f69b891[0]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_977786e4 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[10]),
    .d(al_64a46519[10]),
    .e(al_8a4cc919[10]),
    .o(al_f69b891[10]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_56f23ef6 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[11]),
    .d(al_64a46519[11]),
    .e(al_8a4cc919[11]),
    .o(al_f69b891[11]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_f065b61f (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[12]),
    .d(al_64a46519[12]),
    .e(al_8a4cc919[12]),
    .o(al_f69b891[12]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_9588d51a (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[13]),
    .d(al_64a46519[13]),
    .e(al_8a4cc919[13]),
    .o(al_f69b891[13]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_ab7aed40 (
    .a(al_a9476246[0]),
    .b(al_a9476246[1]),
    .c(al_a9476246[2]),
    .d(al_a9476246[3]),
    .o(al_38ceef8c));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_9cced4f0 (
    .a(al_f55c93aa),
    .b(al_f9514cde),
    .c(al_6127633d),
    .o(al_c92c521a));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*A)"),
    .INIT(32'h00200000))
    al_d2679e6b (
    .a(al_38ceef8c),
    .b(al_452dacc5),
    .c(al_23e59594),
    .d(al_a9476246[4]),
    .e(al_a9476246[5]),
    .o(al_da725511));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_898cab04 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[14]),
    .d(al_64a46519[14]),
    .e(al_8a4cc919[14]),
    .o(al_f69b891[14]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_bc660eb9 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[15]),
    .d(al_64a46519[15]),
    .e(al_8a4cc919[15]),
    .o(al_f69b891[15]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_7a678a82 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[1]),
    .d(al_64a46519[1]),
    .e(al_8a4cc919[1]),
    .o(al_f69b891[1]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_ef6b956d (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[2]),
    .d(al_64a46519[2]),
    .e(al_8a4cc919[2]),
    .o(al_f69b891[2]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_897416a2 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[3]),
    .d(al_64a46519[3]),
    .e(al_8a4cc919[3]),
    .o(al_f69b891[3]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_db600156 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[4]),
    .d(al_64a46519[4]),
    .e(al_8a4cc919[4]),
    .o(al_f69b891[4]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_add210f7 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[5]),
    .d(al_64a46519[5]),
    .e(al_8a4cc919[5]),
    .o(al_f69b891[5]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_5be59503 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[6]),
    .d(al_64a46519[6]),
    .e(al_8a4cc919[6]),
    .o(al_f69b891[6]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_bbf28d5e (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[7]),
    .d(al_64a46519[7]),
    .e(al_8a4cc919[7]),
    .o(al_f69b891[7]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_894f462a (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[8]),
    .d(al_64a46519[8]),
    .e(al_8a4cc919[8]),
    .o(al_f69b891[8]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_5f291270 (
    .a(al_da725511),
    .b(al_c92c521a),
    .c(al_7d74a9c[9]),
    .d(al_64a46519[9]),
    .e(al_8a4cc919[9]),
    .o(al_f69b891[9]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    al_870bfe5f (
    .a(al_520772a3[0]),
    .b(al_452dacc5),
    .c(al_a9476246[0]),
    .o(al_81fd75dc[0]));
  AL_MAP_LUT4 #(
    .EQN("((D@C)*~(B*A))"),
    .INIT(16'h0770))
    al_db462662 (
    .a(al_520772a3[0]),
    .b(al_452dacc5),
    .c(al_a9476246[0]),
    .d(al_a9476246[1]),
    .o(al_81fd75dc[1]));
  AL_MAP_LUT5 #(
    .EQN("((E@(D*C))*~(B*A))"),
    .INIT(32'h07777000))
    al_5b422fed (
    .a(al_520772a3[0]),
    .b(al_452dacc5),
    .c(al_a9476246[0]),
    .d(al_a9476246[1]),
    .e(al_a9476246[2]),
    .o(al_81fd75dc[2]));
  AL_MAP_LUT6 #(
    .EQN("((F@(E*D*C))*~(B*A))"),
    .INIT(64'h0777777770000000))
    al_71f722b6 (
    .a(al_520772a3[0]),
    .b(al_452dacc5),
    .c(al_a9476246[0]),
    .d(al_a9476246[1]),
    .e(al_a9476246[2]),
    .f(al_a9476246[3]),
    .o(al_81fd75dc[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*(D@A))"),
    .INIT(16'h152a))
    al_1560a427 (
    .a(al_38ceef8c),
    .b(al_520772a3[0]),
    .c(al_452dacc5),
    .d(al_a9476246[4]),
    .o(al_81fd75dc[4]));
  AL_MAP_LUT5 #(
    .EQN("(~(C*B)*(E@(D*A)))"),
    .INIT(32'h153f2a00))
    al_341c2875 (
    .a(al_38ceef8c),
    .b(al_520772a3[0]),
    .c(al_452dacc5),
    .d(al_a9476246[4]),
    .e(al_a9476246[5]),
    .o(al_81fd75dc[5]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_fc8756d1 (
    .a(al_64a46519[10]),
    .b(al_64a46519[11]),
    .c(al_64a46519[12]),
    .d(al_64a46519[13]),
    .e(al_64a46519[14]),
    .f(al_64a46519[15]),
    .o(al_de6e30a1));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_3fea8fb9 (
    .a(al_64a46519[4]),
    .b(al_64a46519[5]),
    .c(al_64a46519[6]),
    .d(al_64a46519[7]),
    .e(al_64a46519[8]),
    .f(al_64a46519[9]),
    .o(al_fbe1feab));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_de418e64 (
    .a(al_de6e30a1),
    .b(al_fbe1feab),
    .c(al_64a46519[0]),
    .d(al_64a46519[1]),
    .e(al_64a46519[2]),
    .f(al_64a46519[3]),
    .o(al_240f6a60));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~(C*B)))"),
    .INIT(16'h5540))
    al_418e4c1a (
    .a(al_240f6a60),
    .b(al_520772a3[0]),
    .c(al_9cae7666),
    .d(al_23e59594),
    .o(al_d133c6bf));
  AL_DFF_X al_cb06d5ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d133c6bf),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_23e59594));
  AL_DFF_X al_a46bc817 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[8]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[8]));
  AL_DFF_X al_53f8a1de (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[9]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[9]));
  AL_DFF_X al_9fb175bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[10]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[10]));
  AL_DFF_X al_aa75fa79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[11]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[11]));
  AL_DFF_X al_8771e2a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[12]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[12]));
  AL_DFF_X al_24e21b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[13]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[13]));
  AL_DFF_X al_a5ca1a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[14]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[14]));
  AL_DFF_X al_557c3be (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[15]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[15]));
  AL_DFF_X al_b4338e3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[0]));
  AL_DFF_X al_a7c83e95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[1]));
  AL_DFF_X al_9c534cf0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[2]));
  AL_DFF_X al_b45c7b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[3]));
  AL_DFF_X al_e598d3aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[4]));
  AL_DFF_X al_f5ea35fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[5]));
  AL_DFF_X al_3e5562ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[6]));
  AL_DFF_X al_b6d7dd04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f69b891[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_64a46519[7]));
  AL_DFF_X al_5b369923 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_81fd75dc[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_a9476246[0]));
  AL_DFF_X al_93d5a4ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_81fd75dc[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_a9476246[1]));
  AL_DFF_X al_b951189c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_81fd75dc[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_a9476246[2]));
  AL_DFF_X al_5a2ba8b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_81fd75dc[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_a9476246[3]));
  AL_DFF_X al_6c31930a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_81fd75dc[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_a9476246[4]));
  AL_DFF_X al_cc3fa1f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_81fd75dc[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_a9476246[5]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f7178e0c (
    .a(1'b0),
    .o({al_7c925305,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_54e3a14a (
    .a(al_64a46519[0]),
    .b(1'b1),
    .c(al_7c925305),
    .o({al_41a3eebf,al_8a4cc919[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a60af6ac (
    .a(al_64a46519[1]),
    .b(1'b0),
    .c(al_41a3eebf),
    .o({al_5b5454d7,al_8a4cc919[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_37d17db3 (
    .a(al_64a46519[2]),
    .b(1'b0),
    .c(al_5b5454d7),
    .o({al_a52c4218,al_8a4cc919[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_edfd3c61 (
    .a(al_64a46519[3]),
    .b(1'b0),
    .c(al_a52c4218),
    .o({al_2456cab6,al_8a4cc919[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b46596b3 (
    .a(al_64a46519[4]),
    .b(1'b0),
    .c(al_2456cab6),
    .o({al_c88ff5bc,al_8a4cc919[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_52e33f79 (
    .a(al_64a46519[5]),
    .b(1'b0),
    .c(al_c88ff5bc),
    .o({al_d7c1f764,al_8a4cc919[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_abdcb8ac (
    .a(al_64a46519[6]),
    .b(1'b0),
    .c(al_d7c1f764),
    .o({al_ca164e15,al_8a4cc919[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee2e6904 (
    .a(al_64a46519[7]),
    .b(1'b0),
    .c(al_ca164e15),
    .o({al_6fc51898,al_8a4cc919[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e5328aea (
    .a(al_64a46519[8]),
    .b(1'b0),
    .c(al_6fc51898),
    .o({al_460e3807,al_8a4cc919[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b2e85db7 (
    .a(al_64a46519[9]),
    .b(1'b0),
    .c(al_460e3807),
    .o({al_b1302323,al_8a4cc919[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3f26c8e4 (
    .a(al_64a46519[10]),
    .b(1'b0),
    .c(al_b1302323),
    .o({al_2f1e9be,al_8a4cc919[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6d90b422 (
    .a(al_64a46519[11]),
    .b(1'b0),
    .c(al_2f1e9be),
    .o({al_5617038b,al_8a4cc919[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4885140f (
    .a(al_64a46519[12]),
    .b(1'b0),
    .c(al_5617038b),
    .o({al_7807b4dd,al_8a4cc919[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c3e78511 (
    .a(al_64a46519[13]),
    .b(1'b0),
    .c(al_7807b4dd),
    .o({al_511c2516,al_8a4cc919[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bfed2004 (
    .a(al_64a46519[14]),
    .b(1'b0),
    .c(al_511c2516),
    .o({al_c4a95f07,al_8a4cc919[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4d2549f3 (
    .a(al_64a46519[15]),
    .b(1'b0),
    .c(al_c4a95f07),
    .o({open_n3,al_8a4cc919[15]}));
  AL_DFF_0 al_2f149692 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_47f8fdc1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_58e61c93));
  AL_DFF_0 al_d8a61244 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_58e61c93),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6127633d));
  AL_DFF_X al_17031769 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d1cfb12d),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_retransmit));
  AL_DFF_X al_f89d9cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_stop),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e101ff9a));
  AL_DFF_X al_cb15e0ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_data[0]));
  AL_DFF_X al_fcdb6092 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_data[1]));
  AL_DFF_X al_f42dc070 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_data[2]));
  AL_DFF_X al_4bd6e7f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_data[3]));
  AL_DFF_X al_7b233bcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_data[4]));
  AL_DFF_X al_55c86cd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_data[5]));
  AL_DFF_X al_67b60d02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_data[6]));
  AL_DFF_X al_1c744992 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aeb75558[7]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_data[7]));
  AL_DFF_X al_77bd75a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c01774ad[0]));
  AL_DFF_X al_a02a8bbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c01774ad[1]));
  AL_DFF_X al_b786331b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c01774ad[2]));
  AL_DFF_X al_a8e03bb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c01774ad[3]));
  AL_DFF_X al_7fd7d4d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c01774ad[4]));
  AL_DFF_X al_60b9fdf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c01774ad[5]));
  AL_DFF_X al_cd401401 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c01774ad[6]));
  AL_DFF_X al_8205e2be (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c01774ad[7]));
  AL_DFF_0 al_d74c0e56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_677d00f0[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a7dbaac0));
  AL_DFF_0 al_484ecae6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_a7dbaac0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e495ee45));
  AL_DFF_0 al_8312bf2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_871e6587[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16d49820));
  AL_DFF_0 al_96afda99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_16d49820),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a76fca28));
  AL_DFF_0 al_a3bb56e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_32c99495[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2e8c346));
  AL_DFF_0 al_db66489 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f2e8c346),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715e8e22));
  AL_DFF_0 al_5967fc47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_871e6587[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5a4539df));
  AL_DFF_0 al_df54009d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5a4539df),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_637ddda1));
  AL_DFF_X al_97afb6c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e78cfe9),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_aceaab6b));
  AL_DFF_X al_db761c15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d811499f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d5fb3fbb));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*~D*C*B*A)"),
    .INIT(64'h0000000000800000))
    al_675d4eb7 (
    .a(al_eb34b0be[2]),
    .b(al_eb34b0be[3]),
    .c(al_6ae08f56[0]),
    .d(al_6ae08f56[1]),
    .e(al_6ae08f56[2]),
    .f(al_6ae08f56[3]),
    .o(al_53653f1d));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_d8cc4cd6 (
    .a(al_53653f1d),
    .b(al_eb34b0be[0]),
    .c(al_eb34b0be[1]),
    .o(al_38a4dea8));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_1e740fe1 (
    .a(al_38a4dea8),
    .b(al_2839f3fc),
    .o(al_18862d32));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_31f58f9a (
    .a(al_18862d32),
    .b(al_d5fb3fbb),
    .c(al_fea77e50),
    .o(al_d811499f));
  AL_DFF_X al_7b9d2faa (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fb84638b),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_78920a9b));
  AL_DFF_X al_fab5f976 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_78920a9b),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_6298ef12));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_218696f2 (
    .a(al_124a5ff1),
    .b(al_2d0b2d41),
    .c(al_a533f139),
    .o(al_fb84638b));
  AL_DFF_X al_6f7ce988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rx_vld),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_38ea65b9));
  AL_DFF_X al_870eebc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_38ea65b9),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_124a5ff1));
  AL_DFF_X al_f2022f20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9848ae60),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6842e259));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    al_19d8f933 (
    .a(al_38ea65b9),
    .b(al_124a5ff1),
    .c(al_5c90f2da[0]),
    .d(al_44560df6[1]),
    .o(al_e78cfe9));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(~C*A))"),
    .INIT(16'h00c4))
    al_46e465d9 (
    .a(al_e78cfe9),
    .b(al_124a5ff1),
    .c(al_2d0b2d41),
    .d(al_fea77e50),
    .o(al_9848ae60));
  AL_DFF_X al_69fb2b64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rx_er),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_524c4c86));
  AL_DFF_X al_c0c00683 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_524c4c86),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_2d0b2d41));
  AL_DFF_X al_5268530c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2d0b2d41),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7ca091b));
  AL_DFF_X al_70842859 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7ca091b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e1e36fb));
  AL_DFF_X al_59cf083d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_18862d32),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f4745b25));
  AL_DFF_X al_9e0bb6e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f4745b25),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_a533f139));
  AL_MAP_LUT6 #(
    .EQN("~(~(~C*B)*~(F*~(~E*~D*A)))"),
    .INIT(64'hffffff5d0c0c0c0c))
    al_6be60c7f (
    .a(al_38a4dea8),
    .b(al_38ea65b9),
    .c(al_124a5ff1),
    .d(al_524c4c86),
    .e(al_2d0b2d41),
    .f(al_2839f3fc),
    .o(al_16bdb356));
  AL_DFF_X al_eb5ca101 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_16bdb356),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_2839f3fc));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e1e2945c (
    .a(al_124a5ff1),
    .b(al_5c90f2da[0]),
    .o(al_d19ca65b));
  AL_DFF_X al_ec3423c7 (
    .ar(al_2839f3fc),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d19ca65b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5c90f2da[0]));
  AL_DFF_X al_5c79fc43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[0]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_eb34b0be[0]));
  AL_DFF_X al_88f731f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[1]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_eb34b0be[1]));
  AL_DFF_X al_d2a8a0b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[2]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_eb34b0be[2]));
  AL_DFF_X al_ad44ac82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[3]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_eb34b0be[3]));
  AL_DFF_X al_a61e72ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[4]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_eb34b0be[4]));
  AL_DFF_X al_8b12691f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[5]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_eb34b0be[5]));
  AL_DFF_X al_67a89d51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[6]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_eb34b0be[6]));
  AL_DFF_X al_4e2d8473 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[7]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_eb34b0be[7]));
  AL_DFF_X al_6597d210 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_eb34b0be[0]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_6ae08f56[0]));
  AL_DFF_X al_a6865f08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_eb34b0be[1]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_6ae08f56[1]));
  AL_DFF_X al_5b9e9552 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_eb34b0be[2]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_6ae08f56[2]));
  AL_DFF_X al_e6b4885c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_eb34b0be[3]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_6ae08f56[3]));
  AL_DFF_X al_dba9812f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6ae08f56[0]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f0ba390f[0]));
  AL_DFF_X al_1f3e43eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6ae08f56[1]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f0ba390f[1]));
  AL_DFF_X al_b357ed62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6ae08f56[2]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f0ba390f[2]));
  AL_DFF_X al_1366142b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6ae08f56[3]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f0ba390f[3]));
  AL_DFF_X al_44958aef (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0ba390f[0]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_2fda9ea8[0]));
  AL_DFF_X al_d35aedeb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0ba390f[1]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_2fda9ea8[1]));
  AL_DFF_X al_28678c7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0ba390f[2]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_2fda9ea8[2]));
  AL_DFF_X al_cb7b1f78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0ba390f[3]),
    .en(1'b1),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_2fda9ea8[3]));
  AL_DFF_X al_5c8be4b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(gmii_col),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_22f0d00f));
  AL_DFF_X al_ed609d6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_22f0d00f),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_33156af5));
  AL_DFF_X al_3bb94c0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3daf6177),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_8f006d4e));
  AL_DFF_X al_671c7832 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8f006d4e),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_de5e814a));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'h333305af))
    al_12058c8e (
    .a(al_66d7ef91),
    .b(al_f279ca9c[0]),
    .c(al_be455f81[0]),
    .d(al_be455f81[4]),
    .e(al_44560df6[1]),
    .o(al_fec67178));
  AL_MAP_LUT5 #(
    .EQN("~(~(~C*~B)*~(~E*~(D*~A)))"),
    .INIT(32'h0303abff))
    al_24ad85ae (
    .a(al_b436d586),
    .b(al_197bd181),
    .c(al_fec67178),
    .d(al_8f160d47),
    .e(al_a0ae817c),
    .o(al_3b8f6a2b[0]));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'h333305af))
    al_73c41368 (
    .a(al_66d7ef91),
    .b(al_f279ca9c[1]),
    .c(al_be455f81[1]),
    .d(al_be455f81[5]),
    .e(al_44560df6[1]),
    .o(al_587464d));
  AL_MAP_LUT5 #(
    .EQN("~(~(~C*~B)*~(~E*~(D*~A)))"),
    .INIT(32'h0303abff))
    al_f16cfb8b (
    .a(al_b436d586),
    .b(al_197bd181),
    .c(al_587464d),
    .d(al_8f160d47),
    .e(al_a0ae817c),
    .o(al_3b8f6a2b[1]));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'h333305af))
    al_d49f5cce (
    .a(al_66d7ef91),
    .b(al_f279ca9c[2]),
    .c(al_be455f81[2]),
    .d(al_be455f81[6]),
    .e(al_44560df6[1]),
    .o(al_df75d779));
  AL_MAP_LUT5 #(
    .EQN("~(~(~C*~B)*~(~E*~(D*~A)))"),
    .INIT(32'h0303abff))
    al_8ef72f6f (
    .a(al_b436d586),
    .b(al_197bd181),
    .c(al_df75d779),
    .d(al_8f160d47),
    .e(al_a0ae817c),
    .o(al_3b8f6a2b[2]));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'h333305af))
    al_21804f7d (
    .a(al_66d7ef91),
    .b(al_f279ca9c[3]),
    .c(al_be455f81[3]),
    .d(al_be455f81[7]),
    .e(al_44560df6[1]),
    .o(al_10c967cd));
  AL_MAP_LUT5 #(
    .EQN("~(~(~C*~B)*~(~E*~(D*~A)))"),
    .INIT(32'h0303abff))
    al_ee7c41f6 (
    .a(al_b436d586),
    .b(al_197bd181),
    .c(al_10c967cd),
    .d(al_8f160d47),
    .e(al_a0ae817c),
    .o(al_3b8f6a2b[3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_41e112d8 (
    .a(al_ecabfff7[0]),
    .b(al_ecabfff7[1]),
    .c(al_ecabfff7[2]),
    .d(al_ecabfff7[3]),
    .o(al_8f160d47));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((~E*~D)*~((~C*~B))*~(F)+(~E*~D)*(~C*~B)*~(F)+~((~E*~D))*(~C*~B)*F+(~E*~D)*(~C*~B)*F))"),
    .INIT(64'h5454545455555500))
    al_4312db7c (
    .a(al_f55cb982),
    .b(al_302d0d8b[3]),
    .c(al_302d0d8b[5]),
    .d(al_302d0d8b[7]),
    .e(al_302d0d8b[11]),
    .f(al_44560df6[1]),
    .o(al_197bd181));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~B)*~(~D*~(C*~A)))"),
    .INIT(64'h33bf00af00af00af))
    al_eb0ccdf6 (
    .a(al_b436d586),
    .b(al_197bd181),
    .c(al_8f160d47),
    .d(al_a0ae817c),
    .e(al_f279ca9c[4]),
    .f(al_44560df6[1]),
    .o(al_3b8f6a2b[4]));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~D*~C*~B*A)"),
    .INIT(32'hfffffffd))
    al_b3e9ef7a (
    .a(al_8f160d47),
    .b(al_e08d2b14[0]),
    .c(al_e08d2b14[1]),
    .d(al_e08d2b14[2]),
    .e(al_e08d2b14[3]),
    .o(al_f55cb982));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_a4236068 (
    .a(al_8f006d4e),
    .b(al_de5e814a),
    .c(al_44560df6[1]),
    .o(al_a0ae817c));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h4450))
    al_5e953fe3 (
    .a(al_c5eafaca),
    .b(al_ca7097d4),
    .c(al_48f0356f),
    .d(al_44560df6[1]),
    .o(al_f6f1aa20));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_a8284a41 (
    .a(al_f6f1aa20),
    .b(al_4c8ab20f[0]),
    .c(al_4c8ab20f[1]),
    .d(al_4c8ab20f[2]),
    .e(al_4c8ab20f[3]),
    .o(al_eb5ace4a));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~C*~B))"),
    .INIT(32'haaaaaaa8))
    al_d2e5e616 (
    .a(al_eb5ace4a),
    .b(al_e08d2b14[0]),
    .c(al_e08d2b14[1]),
    .d(al_e08d2b14[2]),
    .e(al_e08d2b14[3]),
    .o(al_b436d586));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(D*A))"),
    .INIT(16'hae0c))
    al_367c77c4 (
    .a(al_1b4e1994),
    .b(al_b436d586),
    .c(al_a0ae817c),
    .d(al_f279ca9c[5]),
    .o(al_3b8f6a2b[5]));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(D*A))"),
    .INIT(16'hae0c))
    al_76c7d5e0 (
    .a(al_1b4e1994),
    .b(al_b436d586),
    .c(al_a0ae817c),
    .d(al_f279ca9c[6]),
    .o(al_3b8f6a2b[6]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_8d87a676 (
    .a(al_8f160d47),
    .b(al_a0ae817c),
    .o(al_a2b6b866));
  AL_MAP_LUT5 #(
    .EQN("(E*~B*~(~A*~(~D*~C)))"),
    .INIT(32'h22230000))
    al_59390778 (
    .a(al_f55cb982),
    .b(al_a2b6b866),
    .c(al_302d0d8b[3]),
    .d(al_302d0d8b[5]),
    .e(al_44560df6[1]),
    .o(al_1b4e1994));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(D*A))"),
    .INIT(16'hae0c))
    al_2f3ac8f9 (
    .a(al_1b4e1994),
    .b(al_b436d586),
    .c(al_a0ae817c),
    .d(al_f279ca9c[7]),
    .o(al_3b8f6a2b[7]));
  AL_DFF_X al_a43e5ec8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_902ad644),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c5eafaca));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e0b3ba5f (
    .a(al_ca7097d4),
    .b(al_48f0356f),
    .c(al_44560df6[1]),
    .o(al_902ad644));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(D*~B*~(~E*~C)))"),
    .INIT(32'hbbaabaaa))
    al_7f0e928f (
    .a(al_b436d586),
    .b(al_197bd181),
    .c(al_8f160d47),
    .d(al_902ad644),
    .e(al_3daf6177),
    .o(al_63772beb));
  AL_DFF_X al_b6ce982a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_63772beb),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d32c67d0));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_e544b61c (
    .a(al_e9410de9),
    .b(al_90130b74),
    .c(al_44560df6[1]),
    .o(al_69a4217a));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~(~E*~C)*~(D*~B)))"),
    .INIT(32'h11001505))
    al_a337f5e3 (
    .a(al_b436d586),
    .b(al_197bd181),
    .c(al_8f160d47),
    .d(al_69a4217a),
    .e(al_3daf6177),
    .o(al_525bf098));
  AL_DFF_X al_4ee35866 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_525bf098),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_31529785));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_86969cb3 (
    .a(al_d1b2b221),
    .b(al_a2b6b866),
    .c(al_ecabfff7[0]),
    .o(al_18a8d68c[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(~C*B)))"),
    .INIT(16'h5104))
    al_e20e761 (
    .a(al_d1b2b221),
    .b(al_a2b6b866),
    .c(al_ecabfff7[0]),
    .d(al_ecabfff7[1]),
    .o(al_18a8d68c[1]));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*D*C*B*~A)"),
    .INIT(64'h0000400000000000))
    al_ac299a8a (
    .a(al_902ad644),
    .b(al_a0ae817c),
    .c(al_69a4217a),
    .d(al_22f0d00f),
    .e(al_33156af5),
    .f(al_32c99495[2]),
    .o(al_d1b2b221));
  AL_MAP_LUT6 #(
    .EQN("((E@(~D*~C*B))*~(F)*~(A)+(E@(~D*~C*B))*F*~(A)+~((E@(~D*~C*B)))*F*A+(E@(~D*~C*B))*F*A)"),
    .INIT(64'hfffbaaae55510004))
    al_4846d725 (
    .a(al_d1b2b221),
    .b(al_a2b6b866),
    .c(al_ecabfff7[0]),
    .d(al_ecabfff7[1]),
    .e(al_ecabfff7[2]),
    .f(al_44560df6[1]),
    .o(al_18a8d68c[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_a09233f0 (
    .a(al_a0ae817c),
    .b(al_ecabfff7[0]),
    .c(al_ecabfff7[1]),
    .d(al_ecabfff7[2]),
    .o(al_713dc35e));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*~B)*~(D)*~(A)+~(C*~B)*D*~(A)+~(~(C*~B))*D*A+~(C*~B)*D*A)"),
    .INIT(16'h10ba))
    al_4b342daf (
    .a(al_d1b2b221),
    .b(al_713dc35e),
    .c(al_ecabfff7[3]),
    .d(al_44560df6[1]),
    .o(al_18a8d68c[3]));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_119ba264 (
    .a(al_b436d586),
    .b(al_aa6b82f0),
    .c(al_e08d2b14[0]),
    .o(al_2ddf456e[0]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(~C*A)))"),
    .INIT(16'h3102))
    al_85875ae6 (
    .a(al_b436d586),
    .b(al_aa6b82f0),
    .c(al_e08d2b14[0]),
    .d(al_e08d2b14[1]),
    .o(al_2ddf456e[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    al_aa05363a (
    .a(al_902ad644),
    .b(al_22f0d00f),
    .c(al_33156af5),
    .d(al_32c99495[2]),
    .o(al_aa6b82f0));
  AL_MAP_LUT6 #(
    .EQN("((E@(~D*~C*A))*~(F)*~(B)+(E@(~D*~C*A))*F*~(B)+~((E@(~D*~C*A)))*F*B+(E@(~D*~C*A))*F*B)"),
    .INIT(64'hfffdccce33310002))
    al_a6310f3c (
    .a(al_b436d586),
    .b(al_aa6b82f0),
    .c(al_e08d2b14[0]),
    .d(al_e08d2b14[1]),
    .e(al_e08d2b14[2]),
    .f(al_44560df6[1]),
    .o(al_2ddf456e[2]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~D*~C*~B*A))"),
    .INIT(32'hfffd0000))
    al_5df6500a (
    .a(al_eb5ace4a),
    .b(al_e08d2b14[0]),
    .c(al_e08d2b14[1]),
    .d(al_e08d2b14[2]),
    .e(al_e08d2b14[3]),
    .o(al_55d8b8f7[3]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'h2e))
    al_e8db2743 (
    .a(al_55d8b8f7[3]),
    .b(al_aa6b82f0),
    .c(al_44560df6[1]),
    .o(al_2ddf456e[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    al_282180da (
    .a(al_66d7ef91),
    .b(al_ca7097d4),
    .c(al_48f0356f),
    .o(al_4462abf6));
  AL_DFF_X al_a992f458 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4462abf6),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_66d7ef91));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    al_221d8acc (
    .a(al_eb5ace4a),
    .b(al_f6f1aa20),
    .c(al_4c8ab20f[0]),
    .o(al_e7fcc128[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*(D@C)))"),
    .INIT(16'h5445))
    al_15078fd0 (
    .a(al_eb5ace4a),
    .b(al_f6f1aa20),
    .c(al_4c8ab20f[0]),
    .d(al_4c8ab20f[1]),
    .o(al_e7fcc128[1]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*(~((~C*~B))*~(D)*~(E)+(~C*~B)*~(D)*~(E)+(~C*~B)*D*~(E)+~((~C*~B))*~(D)*E+(~C*~B)*D*E))"),
    .INIT(32'hfeabfeaa))
    al_c74b9e54 (
    .a(al_f6f1aa20),
    .b(al_4c8ab20f[0]),
    .c(al_4c8ab20f[1]),
    .d(al_4c8ab20f[2]),
    .e(al_4c8ab20f[3]),
    .o(al_e7fcc128[2]));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(~D*~C*~B))*~(F)*~(A)+~(E*~(~D*~C*~B))*F*~(A)+~(~(E*~(~D*~C*~B)))*F*A+~(E*~(~D*~C*~B))*F*A)"),
    .INIT(64'h55540000fffeaaaa))
    al_2438dbaa (
    .a(al_f6f1aa20),
    .b(al_4c8ab20f[0]),
    .c(al_4c8ab20f[1]),
    .d(al_4c8ab20f[2]),
    .e(al_4c8ab20f[3]),
    .f(al_44560df6[1]),
    .o(al_e7fcc128[3]));
  AL_DFF_X al_e96729a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b241735d),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_ca7097d4));
  AL_DFF_X al_530131ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ca7097d4),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_48f0356f));
  AL_DFF_X al_1c729281 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3fc75a33),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e9410de9));
  AL_DFF_X al_ef2b61a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e9410de9),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_90130b74));
  AL_DFF_X al_4acccde1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3b8f6a2b[0]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_42702950[0]));
  AL_DFF_X al_32b3347 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3b8f6a2b[1]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_42702950[1]));
  AL_DFF_X al_90f0886a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3b8f6a2b[2]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_42702950[2]));
  AL_DFF_X al_8bec64fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3b8f6a2b[3]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_42702950[3]));
  AL_DFF_X al_19b3d4fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3b8f6a2b[4]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_42702950[4]));
  AL_DFF_X al_58947518 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3b8f6a2b[5]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_42702950[5]));
  AL_DFF_X al_957729c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3b8f6a2b[6]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_42702950[6]));
  AL_DFF_X al_16f787ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3b8f6a2b[7]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_42702950[7]));
  AL_DFF_X al_1ea4fc90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[7]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[8]));
  AL_DFF_X al_62b8e3f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[8]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[9]));
  AL_DFF_X al_ff69f9fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[9]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[10]));
  AL_DFF_X al_3c99cd6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[10]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[11]));
  AL_DFF_X al_36971d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f55cb982),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[0]));
  AL_DFF_X al_c71ee422 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[0]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[1]));
  AL_DFF_X al_d7ec6e6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[1]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[2]));
  AL_DFF_X al_64fc7775 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[2]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[3]));
  AL_DFF_X al_fc06b7ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[3]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[4]));
  AL_DFF_X al_806bb229 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[4]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[5]));
  AL_DFF_X al_20111736 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[5]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[6]));
  AL_DFF_X al_31060d60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_302d0d8b[6]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_302d0d8b[7]));
  AL_DFF_X al_9242d663 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_18a8d68c[0]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_ecabfff7[0]));
  AL_DFF_X al_9d3ac6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_18a8d68c[1]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_ecabfff7[1]));
  AL_DFF_X al_d94ba700 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_18a8d68c[2]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_ecabfff7[2]));
  AL_DFF_X al_ba3a40da (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_18a8d68c[3]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_ecabfff7[3]));
  AL_DFF_X al_3b6ed44a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ddf456e[0]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e08d2b14[0]));
  AL_DFF_X al_da9c9e05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ddf456e[1]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e08d2b14[1]));
  AL_DFF_X al_644b1170 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ddf456e[2]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e08d2b14[2]));
  AL_DFF_X al_c9dfcf73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ddf456e[3]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e08d2b14[3]));
  AL_DFF_X al_e07c22e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e7fcc128[0]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_4c8ab20f[0]));
  AL_DFF_X al_a8c9bcc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e7fcc128[1]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_4c8ab20f[1]));
  AL_DFF_X al_1031e4ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e7fcc128[2]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_4c8ab20f[2]));
  AL_DFF_X al_1dddfbbc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e7fcc128[3]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_4c8ab20f[3]));
  AL_DFF_X al_1735fb11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f24f9b58[0]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f279ca9c[0]));
  AL_DFF_X al_9c798563 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f24f9b58[1]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f279ca9c[1]));
  AL_DFF_X al_ba043ae0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f24f9b58[2]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f279ca9c[2]));
  AL_DFF_X al_11bfc27d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f24f9b58[3]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f279ca9c[3]));
  AL_DFF_X al_b3fe95a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f24f9b58[4]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f279ca9c[4]));
  AL_DFF_X al_d0a1b832 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f24f9b58[5]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f279ca9c[5]));
  AL_DFF_X al_2b0a12b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f24f9b58[6]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f279ca9c[6]));
  AL_DFF_X al_fef14b83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f24f9b58[7]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f279ca9c[7]));
  AL_DFF_X al_c78f9dce (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f279ca9c[0]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_be455f81[0]));
  AL_DFF_X al_ec22754d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f279ca9c[1]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_be455f81[1]));
  AL_DFF_X al_49d0db82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f279ca9c[2]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_be455f81[2]));
  AL_DFF_X al_c8107279 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f279ca9c[3]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_be455f81[3]));
  AL_DFF_X al_726aad26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f279ca9c[4]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_be455f81[4]));
  AL_DFF_X al_6a293079 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f279ca9c[5]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_be455f81[5]));
  AL_DFF_X al_1b07c22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f279ca9c[6]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_be455f81[6]));
  AL_DFF_X al_4618954a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f279ca9c[7]),
    .en(gmii_tx_clken),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_be455f81[7]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'hccccfa50))
    al_80adf73e (
    .a(al_d5fb3fbb),
    .b(al_eb34b0be[0]),
    .c(al_f0ba390f[0]),
    .d(al_2fda9ea8[0]),
    .e(al_44560df6[1]),
    .o(al_53486c5d[0]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'hccccfa50))
    al_53245b9d (
    .a(al_d5fb3fbb),
    .b(al_eb34b0be[1]),
    .c(al_f0ba390f[1]),
    .d(al_2fda9ea8[1]),
    .e(al_44560df6[1]),
    .o(al_53486c5d[1]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'hccccfa50))
    al_f8969dbf (
    .a(al_d5fb3fbb),
    .b(al_eb34b0be[2]),
    .c(al_f0ba390f[2]),
    .d(al_2fda9ea8[2]),
    .e(al_44560df6[1]),
    .o(al_53486c5d[2]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'hccccfa50))
    al_d475055b (
    .a(al_d5fb3fbb),
    .b(al_eb34b0be[3]),
    .c(al_f0ba390f[3]),
    .d(al_2fda9ea8[3]),
    .e(al_44560df6[1]),
    .o(al_53486c5d[3]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'hccccfa50))
    al_b0092c (
    .a(al_d5fb3fbb),
    .b(al_eb34b0be[4]),
    .c(al_6ae08f56[0]),
    .d(al_f0ba390f[0]),
    .e(al_44560df6[1]),
    .o(al_53486c5d[4]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'hccccfa50))
    al_ff163a8e (
    .a(al_d5fb3fbb),
    .b(al_eb34b0be[5]),
    .c(al_6ae08f56[1]),
    .d(al_f0ba390f[1]),
    .e(al_44560df6[1]),
    .o(al_53486c5d[5]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'hccccfa50))
    al_57479263 (
    .a(al_d5fb3fbb),
    .b(al_eb34b0be[6]),
    .c(al_6ae08f56[2]),
    .d(al_f0ba390f[2]),
    .e(al_44560df6[1]),
    .o(al_53486c5d[6]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(B)*~(E)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*~(E)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*B*E+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*B*E)"),
    .INIT(32'hccccfa50))
    al_4f56308e (
    .a(al_d5fb3fbb),
    .b(al_eb34b0be[7]),
    .c(al_6ae08f56[3]),
    .d(al_f0ba390f[3]),
    .e(al_44560df6[1]),
    .o(al_53486c5d[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_51f0ef02 (
    .a(al_38ea65b9),
    .b(al_6842e259),
    .c(al_44560df6[1]),
    .o(al_16302c3d));
  AL_MAP_LUT5 #(
    .EQN("(~D*~A*~(~E*C*B))"),
    .INIT(32'h00550015))
    al_a1b8d346 (
    .a(al_6298ef12),
    .b(al_124a5ff1),
    .c(al_2d0b2d41),
    .d(al_7ca091b),
    .e(al_a533f139),
    .o(al_44dddc1d));
  AL_MAP_LUT5 #(
    .EQN("(~(A*~(D*B))*~(C)*~(E)+~(A*~(D*B))*C*~(E)+~(~(A*~(D*B)))*C*E+~(A*~(D*B))*C*E)"),
    .INIT(32'hf0f0dd55))
    al_6b5536d3 (
    .a(al_44dddc1d),
    .b(al_d5fb3fbb),
    .c(al_524c4c86),
    .d(al_e1e36fb),
    .e(al_44560df6[1]),
    .o(al_60057698));
  AL_DFF_X al_5db3623c (
    .ar(1'b0),
    .as(reset),
    .clk(s_axi_aclk),
    .d(1'b0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_760b1195));
  AL_DFF_X al_8d0e0c7a (
    .ar(1'b0),
    .as(reset),
    .clk(s_axi_aclk),
    .d(al_760b1195),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22e99ffa));
  AL_DFF_0 al_52144a1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_22e99ffa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b936a4eb));
  AL_DFF_1 al_73ca1626 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_30591f5d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16296d60));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_d0b6cad5 (
    .a(al_22e99ffa),
    .b(al_b936a4eb),
    .o(al_30591f5d));
  AL_DFF_0 al_9a5de81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_fb466fd8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86bf0006));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*(D@A))"),
    .INIT(16'h0102))
    al_5542428e (
    .a(al_c7821d7e),
    .b(al_46dd4bfb),
    .c(al_16296d60),
    .d(al_86bf0006),
    .o(al_fb466fd8));
  AL_MAP_LUT5 #(
    .EQN("~(~(~(E*~D)*B)*~(C*A))"),
    .INIT(32'heca0ecec))
    al_980921ee (
    .a(al_ec112ad9),
    .b(al_1ff3d4e5),
    .c(al_7de51101[0]),
    .d(al_60f51d47),
    .e(al_9439ddc),
    .o(al_68cc6b50));
  AL_DFF_0 al_a70e95db (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_68cc6b50),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_1ff3d4e5));
  AL_DFF_0 al_dc222263 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_5d24a167),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a60f8a1f[2]));
  AL_DFF_0 al_d52b0718 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_d4b6c586),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a60f8a1f[3]));
  AL_DFF_0 al_160a1dbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_240a1ace),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a60f8a1f[4]));
  AL_DFF_0 al_7f71e7b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_27fc47ee),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a60f8a1f[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_94bcd7df (
    .a(al_a60f8a1f[1]),
    .b(al_a60f8a1f[2]),
    .c(al_a60f8a1f[3]),
    .d(al_3f753490[1]),
    .e(al_3f753490[2]),
    .f(al_3f753490[3]),
    .o(al_d38bd427));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_26580192 (
    .a(al_a60f8a1f[0]),
    .b(al_a60f8a1f[4]),
    .c(al_a60f8a1f[5]),
    .d(al_3f753490[0]),
    .e(al_3f753490[4]),
    .f(al_3f753490[5]),
    .o(al_ffb977ef));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_bde6adda (
    .a(al_d38bd427),
    .b(al_ffb977ef),
    .o(al_c7821d7e));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_f4dcea2d (
    .a(al_c7821d7e),
    .b(al_16296d60),
    .o(al_6fbcf05d));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_f8963393 (
    .a(al_6fbcf05d),
    .b(al_a60f8a1f[0]),
    .o(al_c5d247c0));
  AL_MAP_LUT6 #(
    .EQN("(A*(F@(E*D*C*B)))"),
    .INIT(64'h2aaaaaaa80000000))
    al_3607bff4 (
    .a(al_6fbcf05d),
    .b(al_a60f8a1f[0]),
    .c(al_a60f8a1f[1]),
    .d(al_a60f8a1f[2]),
    .e(al_a60f8a1f[3]),
    .f(al_a60f8a1f[4]),
    .o(al_240a1ace));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    al_925b37b4 (
    .a(al_6fbcf05d),
    .b(al_a60f8a1f[0]),
    .c(al_a60f8a1f[1]),
    .o(al_b3b873e8));
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(C*B)))"),
    .INIT(16'h2a80))
    al_6372a70 (
    .a(al_6fbcf05d),
    .b(al_a60f8a1f[0]),
    .c(al_a60f8a1f[1]),
    .d(al_a60f8a1f[2]),
    .o(al_5d24a167));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@(D*C*B)))"),
    .INIT(32'h2aaa8000))
    al_33bea76a (
    .a(al_6fbcf05d),
    .b(al_a60f8a1f[0]),
    .c(al_a60f8a1f[1]),
    .d(al_a60f8a1f[2]),
    .e(al_a60f8a1f[3]),
    .o(al_d4b6c586));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_8819d082 (
    .a(al_a60f8a1f[0]),
    .b(al_a60f8a1f[1]),
    .c(al_a60f8a1f[2]),
    .d(al_a60f8a1f[3]),
    .e(al_a60f8a1f[4]),
    .f(al_a60f8a1f[5]),
    .o(al_c364719f[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_1b670496 (
    .a(al_6fbcf05d),
    .b(al_c364719f[5]),
    .o(al_27fc47ee));
  AL_DFF_0 al_4ebd2d81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_c5d247c0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a60f8a1f[0]));
  AL_DFF_0 al_63f0a73b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_b3b873e8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a60f8a1f[1]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_c10535fe (
    .a(al_665205be),
    .b(s_axi_araddr[0]),
    .c(s_axi_rvalid),
    .d(al_eb5eeaf9[0]),
    .o(al_6f6e3b4e[0]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_19cd7f03 (
    .a(al_665205be),
    .b(s_axi_araddr[1]),
    .c(s_axi_rvalid),
    .d(al_eb5eeaf9[1]),
    .o(al_6f6e3b4e[1]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_495a00d7 (
    .a(al_665205be),
    .b(s_axi_araddr[2]),
    .c(s_axi_rvalid),
    .d(al_eb5eeaf9[2]),
    .o(al_6f6e3b4e[2]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_792e4cfe (
    .a(al_665205be),
    .b(s_axi_araddr[3]),
    .c(s_axi_rvalid),
    .d(al_eb5eeaf9[3]),
    .o(al_6f6e3b4e[3]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_ef343c6f (
    .a(al_665205be),
    .b(s_axi_araddr[4]),
    .c(s_axi_rvalid),
    .d(al_eb5eeaf9[4]),
    .o(al_6f6e3b4e[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_82fd4188 (
    .a(s_axi_arvalid),
    .b(s_axi_arready),
    .o(al_665205be));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_629018c3 (
    .a(al_665205be),
    .b(s_axi_araddr[5]),
    .c(s_axi_rvalid),
    .d(al_eb5eeaf9[5]),
    .o(al_6f6e3b4e[5]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_49640f1a (
    .a(al_665205be),
    .b(s_axi_araddr[6]),
    .c(s_axi_rvalid),
    .d(al_eb5eeaf9[6]),
    .o(al_6f6e3b4e[6]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_3ff5abec (
    .a(al_665205be),
    .b(s_axi_araddr[7]),
    .c(s_axi_rvalid),
    .d(al_eb5eeaf9[7]),
    .o(al_6f6e3b4e[7]));
  AL_DFF_0 al_c5198d4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_665205be),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(s_axi_arready));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_e20ff929 (
    .a(al_450a8cba),
    .b(s_axi_awaddr[0]),
    .c(s_axi_bvalid),
    .d(al_60c7c349[0]),
    .o(al_dbc70e2f[0]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_72d19c8e (
    .a(al_450a8cba),
    .b(s_axi_awaddr[1]),
    .c(s_axi_bvalid),
    .d(al_60c7c349[1]),
    .o(al_dbc70e2f[1]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_b26c8fda (
    .a(al_450a8cba),
    .b(s_axi_awaddr[2]),
    .c(s_axi_bvalid),
    .d(al_60c7c349[2]),
    .o(al_dbc70e2f[2]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_b7bb521f (
    .a(al_450a8cba),
    .b(s_axi_awaddr[3]),
    .c(s_axi_bvalid),
    .d(al_60c7c349[3]),
    .o(al_dbc70e2f[3]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_9b21d63a (
    .a(al_450a8cba),
    .b(s_axi_awaddr[4]),
    .c(s_axi_bvalid),
    .d(al_60c7c349[4]),
    .o(al_dbc70e2f[4]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_28be2346 (
    .a(s_axi_awvalid),
    .b(s_axi_wvalid),
    .c(s_axi_awready),
    .o(al_450a8cba));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_640764ee (
    .a(al_450a8cba),
    .b(s_axi_awaddr[5]),
    .c(s_axi_bvalid),
    .d(al_60c7c349[5]),
    .o(al_dbc70e2f[5]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_c2c46301 (
    .a(al_450a8cba),
    .b(s_axi_awaddr[6]),
    .c(s_axi_bvalid),
    .d(al_60c7c349[6]),
    .o(al_dbc70e2f[6]));
  AL_MAP_LUT4 #(
    .EQN("((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .INIT(16'h8d88))
    al_9686aaca (
    .a(al_450a8cba),
    .b(s_axi_awaddr[7]),
    .c(s_axi_bvalid),
    .d(al_60c7c349[7]),
    .o(al_dbc70e2f[7]));
  AL_DFF_0 al_96c2e513 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_450a8cba),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(s_axi_awready));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~((F*~E))+~(A)*B*C*~(D)*~((F*~E))+~(A)*~(B)*~(C)*D*~((F*~E))+A*~(B)*~(C)*D*~((F*~E))+~(A)*B*~(C)*D*~((F*~E))+A*B*~(C)*D*~((F*~E))+A*~(B)*~(C)*~(D)*(F*~E)+~(A)*B*~(C)*~(D)*(F*~E)+A*B*~(C)*~(D)*(F*~E)+A*~(B)*C*~(D)*(F*~E)+~(A)*B*C*~(D)*(F*~E)+A*B*C*~(D)*(F*~E)+~(A)*~(B)*~(C)*D*(F*~E)+A*~(B)*~(C)*D*(F*~E)+~(A)*B*~(C)*D*(F*~E)+A*B*~(C)*D*(F*~E)+A*~(B)*C*D*(F*~E)+A*B*C*D*(F*~E))"),
    .INIT(64'h0f44afee0f440f44))
    al_33e28d2a (
    .a(al_b37ae739),
    .b(al_26874532),
    .c(s_axi_bready),
    .d(s_axi_bvalid),
    .e(al_60f51d47),
    .f(al_9439ddc),
    .o(al_b14c08d7));
  AL_DFF_0 al_78939d81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_b14c08d7),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(s_axi_bvalid));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_df9d9de4 (
    .a(s_axi_arvalid),
    .b(s_axi_arready),
    .c(s_axi_rvalid),
    .o(al_5a17606d));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*A)"),
    .INIT(32'h00200000))
    al_47299776 (
    .a(al_8b7519f2),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_eb5eeaf9[6]),
    .e(al_eb5eeaf9[7]),
    .o(al_14c1bc93));
  AL_MAP_LUT6 #(
    .EQN("~(~(D*~C)*~(B*~((F*~E))*~(A)+B*(F*~E)*~(A)+~(B)*(F*~E)*A+B*(F*~E)*A))"),
    .INIT(64'h4f44efee4f444f44))
    al_dab2bc8a (
    .a(al_14c1bc93),
    .b(al_5a17606d),
    .c(s_axi_rready),
    .d(s_axi_rvalid),
    .e(al_60f51d47),
    .f(al_9439ddc),
    .o(al_9cc4302));
  AL_DFF_0 al_600e49c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9cc4302),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(s_axi_rvalid));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*A)"),
    .INIT(32'h02000000))
    al_d28d652 (
    .a(al_9daabc69),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_cee59967));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    al_76948249 (
    .a(al_9daabc69),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_9ec235f9));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_e6e76a0e (
    .a(al_9ec235f9),
    .b(s_axi_wdata[0]),
    .o(al_8ba03385));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_2937481c (
    .a(al_9daabc69),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_8b9cbde3));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_7f50c5e0 (
    .a(al_8b9cbde3),
    .b(s_axi_wdata[0]),
    .o(al_76f4f274));
  AL_DFF_1 al_118ac2c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_d7515c44),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4ebb1964));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    al_f269a2ba (
    .a(al_9daabc69),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_a4aaca2e));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hfdf8))
    al_fcef3bac (
    .a(al_a4aaca2e),
    .b(s_axi_wdata[0]),
    .c(al_16296d60),
    .d(al_4ebb1964),
    .o(al_d7515c44));
  AL_DFF_0 al_4615909b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6f6e3b4e[0]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_eb5eeaf9[0]));
  AL_DFF_0 al_fbcc55e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6f6e3b4e[1]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_eb5eeaf9[1]));
  AL_DFF_0 al_bb88f752 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6f6e3b4e[2]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_eb5eeaf9[2]));
  AL_DFF_0 al_90768ee6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6f6e3b4e[3]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_eb5eeaf9[3]));
  AL_DFF_0 al_6969d743 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6f6e3b4e[4]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_eb5eeaf9[4]));
  AL_DFF_0 al_952f1fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6f6e3b4e[5]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_eb5eeaf9[5]));
  AL_DFF_0 al_57bfbe5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6f6e3b4e[6]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_eb5eeaf9[6]));
  AL_DFF_0 al_51544c40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6f6e3b4e[7]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_eb5eeaf9[7]));
  AL_DFF_0 al_7362b601 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[0]));
  AL_DFF_0 al_2a5c6022 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[1]));
  AL_DFF_0 al_311a11a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[2]));
  AL_DFF_0 al_2e762209 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[3]));
  AL_DFF_0 al_aeca3b57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[4]));
  AL_DFF_0 al_4cae96e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[5]));
  AL_DFF_0 al_c11e6adc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[6]));
  AL_DFF_0 al_732f6f20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[7]));
  AL_DFF_0 al_c7b40d5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[8]));
  AL_DFF_0 al_34adc6b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[9]));
  AL_DFF_0 al_9cf2cf8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[10]));
  AL_DFF_0 al_e62e5a2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[11]));
  AL_DFF_0 al_8661cdc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[12]));
  AL_DFF_0 al_a47b3a12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[13]));
  AL_DFF_0 al_3c68b5b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[14]));
  AL_DFF_0 al_29bda30d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1062ede0[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3c2ad2a[15]));
  AL_DFF_0 al_50ff046a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_8ba03385),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_677d00f0[0]));
  AL_DFF_0 al_5beee436 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[2]));
  AL_DFF_0 al_fb513d68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[3]));
  AL_DFF_0 al_6b9b2042 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[4]));
  AL_DFF_0 al_664fc30f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[5]));
  AL_DFF_0 al_b3e837be (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[6]));
  AL_DFF_0 al_922d492b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[7]));
  AL_DFF_0 al_195d5895 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[8]));
  AL_DFF_0 al_e76a05d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[9]));
  AL_DFF_0 al_d44aac2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[10]));
  AL_DFF_0 al_48e389 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[11]));
  AL_DFF_0 al_d7e493a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[12]));
  AL_DFF_0 al_92d811e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[13]));
  AL_DFF_0 al_4ba8c4c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[14]));
  AL_DFF_0 al_f78faae9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[15]));
  AL_DFF_0 al_eaa2bc40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[16]));
  AL_DFF_0 al_22777be4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[17]));
  AL_DFF_0 al_e2cb1428 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[18]));
  AL_DFF_0 al_d361d63e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[19]));
  AL_DFF_0 al_e76c6506 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[20]));
  AL_DFF_0 al_729ad83a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[21]));
  AL_DFF_0 al_87a1356e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[22]));
  AL_DFF_0 al_2342f439 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[23]));
  AL_DFF_0 al_faa8f23c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[24]));
  AL_DFF_0 al_12488ae5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[25]));
  AL_DFF_0 al_1a66a7ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[26]));
  AL_DFF_0 al_2ab41aaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[27]));
  AL_DFF_0 al_2e923e90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[28]));
  AL_DFF_0 al_4450403e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[29]));
  AL_DFF_0 al_5587d69f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[30]));
  AL_DFF_0 al_9c6bb2b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_9ec235f9),
    .sr(al_655c284a),
    .ss(1'b0),
    .q(al_677d00f0[31]));
  AL_DFF_1 al_dfdca557 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_9ec235f9),
    .sr(1'b0),
    .ss(al_655c284a),
    .q(al_677d00f0[1]));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    al_b292d81f (
    .a(al_9daabc69),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_a360ff8));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_cd66c72d (
    .a(al_a360ff8),
    .b(s_axi_wdata[0]),
    .c(al_44560df6[0]),
    .o(al_39b879bd));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_de530f92 (
    .a(al_a360ff8),
    .b(s_axi_wdata[1]),
    .c(al_44560df6[1]),
    .o(al_dd95f235));
  AL_DFF_0 al_ae324853 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_39b879bd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44560df6[0]));
  AL_DFF_0 al_29a7f0f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dd95f235),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44560df6[1]));
  AL_DFF_0 al_689dc403 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_76f4f274),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_32c99495[0]));
  AL_DFF_0 al_88bd299 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[2]));
  AL_DFF_0 al_db54786e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[3]));
  AL_DFF_0 al_bf073915 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[4]));
  AL_DFF_0 al_f28d9795 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[5]));
  AL_DFF_0 al_5d7fba36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[6]));
  AL_DFF_0 al_66c4dde7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[7]));
  AL_DFF_0 al_2fef98ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[8]));
  AL_DFF_0 al_9c77a249 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[9]));
  AL_DFF_0 al_4b59b105 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[10]));
  AL_DFF_0 al_97a98f4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[11]));
  AL_DFF_0 al_d53e1319 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[12]));
  AL_DFF_0 al_9cda5a4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[13]));
  AL_DFF_0 al_137b8505 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[14]));
  AL_DFF_0 al_b0c2f41e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[15]));
  AL_DFF_0 al_49a8ff52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[16]));
  AL_DFF_0 al_42dfab10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[17]));
  AL_DFF_0 al_d59cea5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[18]));
  AL_DFF_0 al_b0025fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[19]));
  AL_DFF_0 al_a0a97ad1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[20]));
  AL_DFF_0 al_28081d7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[21]));
  AL_DFF_0 al_a36f0c56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[22]));
  AL_DFF_0 al_f7d2b42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[23]));
  AL_DFF_0 al_736b711d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[24]));
  AL_DFF_0 al_714d53eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[25]));
  AL_DFF_0 al_aa99d7e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[26]));
  AL_DFF_0 al_f40a04d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[27]));
  AL_DFF_0 al_1264e279 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[28]));
  AL_DFF_0 al_471df679 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[29]));
  AL_DFF_0 al_a5624a4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[30]));
  AL_DFF_0 al_e83d3d1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_8b9cbde3),
    .sr(al_7fda1410),
    .ss(1'b0),
    .q(al_32c99495[31]));
  AL_DFF_1 al_6f9c08c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_8b9cbde3),
    .sr(1'b0),
    .ss(al_7fda1410),
    .q(al_32c99495[1]));
  AL_DFF_0 al_634483ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dbc70e2f[0]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_60c7c349[0]));
  AL_DFF_0 al_4b42d9bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dbc70e2f[1]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_60c7c349[1]));
  AL_DFF_0 al_4875a90d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dbc70e2f[2]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_60c7c349[2]));
  AL_DFF_0 al_501a3cda (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dbc70e2f[3]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_60c7c349[3]));
  AL_DFF_0 al_7635fbfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dbc70e2f[4]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_60c7c349[4]));
  AL_DFF_0 al_db9e2660 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dbc70e2f[5]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_60c7c349[5]));
  AL_DFF_0 al_1216882a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dbc70e2f[6]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_60c7c349[6]));
  AL_DFF_0 al_7eeca957 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dbc70e2f[7]),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_60c7c349[7]));
  AL_DFF_0 al_44b33054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[0]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[0]));
  AL_DFF_0 al_969d84c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[1]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[1]));
  AL_DFF_0 al_c494eb49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[2]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[2]));
  AL_DFF_0 al_6da9a679 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[3]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[3]));
  AL_DFF_0 al_5394d4fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[4]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[4]));
  AL_DFF_0 al_426ae04f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[5]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[5]));
  AL_DFF_0 al_bbea675 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[6]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[6]));
  AL_DFF_0 al_c807437d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[7]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[7]));
  AL_DFF_0 al_2defb7e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[8]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[8]));
  AL_DFF_0 al_a62d7e38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[9]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[9]));
  AL_DFF_0 al_8defd1f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[10]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[10]));
  AL_DFF_0 al_9aea2046 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[11]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[11]));
  AL_DFF_0 al_235ba8ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[12]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[12]));
  AL_DFF_0 al_7bf91c73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[13]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[13]));
  AL_DFF_0 al_1f632a0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[14]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[14]));
  AL_DFF_0 al_597cb1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[15]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[15]));
  AL_DFF_0 al_8a226fb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[16]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[16]));
  AL_DFF_0 al_48e3f5d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[17]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[17]));
  AL_DFF_0 al_cac6a869 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[18]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[18]));
  AL_DFF_0 al_53acc617 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[19]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[19]));
  AL_DFF_0 al_5fd3c3b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[20]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[20]));
  AL_DFF_0 al_d82ccb65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[21]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[21]));
  AL_DFF_0 al_c702e201 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[22]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[22]));
  AL_DFF_0 al_c6e434a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[23]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[23]));
  AL_DFF_0 al_b334c7dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[24]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[24]));
  AL_DFF_0 al_d0a29499 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[25]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[25]));
  AL_DFF_0 al_5d585822 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[26]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[26]));
  AL_DFF_0 al_7bc1ecd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[27]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[27]));
  AL_DFF_0 al_a22ed29c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[28]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[28]));
  AL_DFF_0 al_7448121a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[29]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[29]));
  AL_DFF_0 al_888a11a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[30]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[30]));
  AL_DFF_0 al_8773a79e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4197a0a2[31]),
    .en(al_5a17606d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_fa4d6e00[31]));
  AL_DFF_1 al_75570f24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_41fb49d4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_871e6587[0]));
  AL_DFF_1 al_e2006fc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_937f8e6e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_871e6587[1]));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*~B*A)"),
    .INIT(32'h00002000))
    al_c61a703c (
    .a(al_9daabc69),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_31ede2e2));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hfdf8))
    al_5ddc03fa (
    .a(al_31ede2e2),
    .b(s_axi_wdata[0]),
    .c(al_16296d60),
    .d(al_871e6587[0]),
    .o(al_41fb49d4));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hfdf8))
    al_f7c4f0f1 (
    .a(al_31ede2e2),
    .b(s_axi_wdata[1]),
    .c(al_16296d60),
    .d(al_871e6587[1]),
    .o(al_937f8e6e));
  AL_DFF_0 al_7b090315 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_f6f8b1fe),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3f753490[1]));
  AL_DFF_0 al_27f6d8d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_fcdf9700),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3f753490[2]));
  AL_DFF_0 al_800de96f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_919f4410),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3f753490[3]));
  AL_DFF_0 al_c07e0b51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_8a13cd79),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3f753490[4]));
  AL_DFF_0 al_7800c426 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_38bb9e5e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3f753490[5]));
  AL_DFF_1 al_766a6a8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_efdfec25),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3f753490[6]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    al_ffc34994 (
    .a(al_9daabc69),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_c291f47d));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_cf966166 (
    .a(al_c291f47d),
    .b(s_axi_wdata[5]),
    .c(al_16296d60),
    .d(al_3f753490[5]),
    .o(al_38bb9e5e));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_8c8ec99e (
    .a(al_c291f47d),
    .b(s_axi_wdata[4]),
    .c(al_16296d60),
    .d(al_3f753490[4]),
    .o(al_8a13cd79));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_5abcb9c1 (
    .a(al_c291f47d),
    .b(s_axi_wdata[0]),
    .c(al_16296d60),
    .d(al_3f753490[0]),
    .o(al_d1b5a8f4));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_16d1ed12 (
    .a(al_c291f47d),
    .b(s_axi_wdata[1]),
    .c(al_16296d60),
    .d(al_3f753490[1]),
    .o(al_f6f8b1fe));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_c7ad5db0 (
    .a(al_c291f47d),
    .b(s_axi_wdata[2]),
    .c(al_16296d60),
    .d(al_3f753490[2]),
    .o(al_fcdf9700));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_e765aab0 (
    .a(al_c291f47d),
    .b(s_axi_wdata[3]),
    .c(al_16296d60),
    .d(al_3f753490[3]),
    .o(al_919f4410));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hfdf8))
    al_9db045d2 (
    .a(al_c291f47d),
    .b(s_axi_wdata[6]),
    .c(al_16296d60),
    .d(al_3f753490[6]),
    .o(al_efdfec25));
  AL_DFF_0 al_f9797478 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_d1b5a8f4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3f753490[0]));
  AL_DFF_0 al_a6e2f104 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_a2d51717),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7de51101[0]));
  AL_DFF_0 al_1cfef376 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[1]));
  AL_DFF_0 al_9a1d5aab (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[2]));
  AL_DFF_0 al_b68a114d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[3]));
  AL_DFF_0 al_76128b47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[4]));
  AL_DFF_0 al_bf560b85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[5]));
  AL_DFF_0 al_9506fb2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[6]));
  AL_DFF_0 al_76c5f961 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[7]));
  AL_DFF_0 al_b22434b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[8]));
  AL_DFF_0 al_86174c97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[9]));
  AL_DFF_0 al_ac4166c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[10]));
  AL_DFF_0 al_473ee077 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[11]));
  AL_DFF_0 al_8eba7765 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_b8f3be80),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_7de51101[12]));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000100000000))
    al_93089e94 (
    .a(al_60c7c349[0]),
    .b(al_60c7c349[1]),
    .c(al_60c7c349[2]),
    .d(al_60c7c349[3]),
    .e(al_60c7c349[4]),
    .f(al_60c7c349[5]),
    .o(al_594ca757));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_ab5a9d20 (
    .a(al_594ca757),
    .b(al_60c7c349[6]),
    .c(al_60c7c349[7]),
    .o(al_b37ae739));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_536c9307 (
    .a(al_b37ae739),
    .b(al_26874532),
    .o(al_b8f3be80));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_23cfdc38 (
    .a(al_b8f3be80),
    .b(s_axi_wdata[0]),
    .c(al_16296d60),
    .d(al_7de51101[0]),
    .o(al_a2d51717));
  AL_DFF_0 al_52f340c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[0]));
  AL_DFF_0 al_90c795b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[1]));
  AL_DFF_0 al_5c6f314a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[2]));
  AL_DFF_0 al_921efae (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[3]));
  AL_DFF_0 al_92d190a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[4]));
  AL_DFF_0 al_1e32f878 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[5]));
  AL_DFF_0 al_9343ea40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[6]));
  AL_DFF_0 al_938332d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[7]));
  AL_DFF_0 al_8c01f334 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[8]));
  AL_DFF_0 al_13c48284 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[9]));
  AL_DFF_0 al_7b74884d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[10]));
  AL_DFF_0 al_4edd5a06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[11]));
  AL_DFF_0 al_475c13ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[12]));
  AL_DFF_0 al_2145b5e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[13]));
  AL_DFF_0 al_7dbd33fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[14]));
  AL_DFF_0 al_807ce766 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_cee59967),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3cae1837[15]));
  AL_DFF_0 al_1762af29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[0]));
  AL_DFF_0 al_e746863a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[1]));
  AL_DFF_0 al_89a74810 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[2]));
  AL_DFF_0 al_da7cd5de (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[3]));
  AL_DFF_0 al_a31fb831 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[4]));
  AL_DFF_0 al_921a97e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[5]));
  AL_DFF_0 al_a93c86dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[6]));
  AL_DFF_0 al_5c8f2fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[7]));
  AL_DFF_0 al_ba7e5ce9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[8]));
  AL_DFF_0 al_3d17a1f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[9]));
  AL_DFF_0 al_19a39180 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[10]));
  AL_DFF_0 al_d8c1d97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[11]));
  AL_DFF_0 al_6b01db35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[12]));
  AL_DFF_0 al_5da9bead (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[13]));
  AL_DFF_0 al_95201da5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[14]));
  AL_DFF_0 al_561d2c94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[15]));
  AL_DFF_0 al_929cba28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[16]));
  AL_DFF_0 al_c9fb2a2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[17]));
  AL_DFF_0 al_a0502821 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[18]));
  AL_DFF_0 al_9a8a6c5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[19]));
  AL_DFF_0 al_8ec396b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[20]));
  AL_DFF_0 al_2e696729 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[21]));
  AL_DFF_0 al_8b40fc20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[22]));
  AL_DFF_0 al_49219729 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[23]));
  AL_DFF_0 al_20074d5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[24]));
  AL_DFF_0 al_2a8e7d07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[25]));
  AL_DFF_0 al_1eb74af4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[26]));
  AL_DFF_0 al_2866d6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[27]));
  AL_DFF_0 al_356ab9df (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[28]));
  AL_DFF_0 al_d69d7beb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[29]));
  AL_DFF_0 al_ab97f297 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[30]));
  AL_DFF_0 al_54ef975c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ae69e57d[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_42381c95[31]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h4567cdef))
    al_52c12661 (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[7]),
    .c(al_677d00f0[0]),
    .d(al_42381c95[0]),
    .e(al_1cb63986[0]),
    .o(al_bdab8dd4));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C))*~(D)+~A*(E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C)*~(D)+~(~A)*(E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C)*D+~A*(E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C)*D)"),
    .INIT(32'h30aa3faa))
    al_6e6aaff1 (
    .a(al_bdab8dd4),
    .b(al_4ebb1964),
    .c(al_eb5eeaf9[4]),
    .d(al_eb5eeaf9[6]),
    .e(al_871e6587[0]),
    .o(al_2156b30e));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_30dd8954 (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[0]),
    .c(al_44560df6[0]),
    .o(al_a100d2c5[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfbf8cbc83b380b08))
    al_b169302b (
    .a(al_a100d2c5[0]),
    .b(al_eb5eeaf9[6]),
    .c(al_eb5eeaf9[7]),
    .d(al_32c99495[0]),
    .e(al_3f753490[0]),
    .f(al_3cae1837[0]),
    .o(al_55bc11eb));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .INIT(16'h44c0))
    al_1bbf0630 (
    .a(al_2156b30e),
    .b(al_e2aa4ae4),
    .c(al_55bc11eb),
    .d(al_eb5eeaf9[5]),
    .o(al_4197a0a2[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_3043a861 (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[10]),
    .o(al_a100d2c5[10]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hc3dff3dfcfdfffdf))
    al_c4618f88 (
    .a(al_a100d2c5[10]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .e(al_3cae1837[10]),
    .f(al_1cb63986[10]),
    .o(al_72a9a166));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*~(B)+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(B)+~(D)*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B)"),
    .INIT(32'h04378cbf))
    al_fc967549 (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_677d00f0[10]),
    .d(al_32c99495[10]),
    .e(al_42381c95[10]),
    .o(al_b58b5a6));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(~D*A))"),
    .INIT(16'h0cae))
    al_798fa457 (
    .a(al_f4b9a391),
    .b(al_e2aa4ae4),
    .c(al_72a9a166),
    .d(al_b58b5a6),
    .o(al_4197a0a2[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b50feba6 (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[11]),
    .o(al_a100d2c5[11]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hc3dff3dfcfdfffdf))
    al_b059a668 (
    .a(al_a100d2c5[11]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .e(al_3cae1837[11]),
    .f(al_1cb63986[11]),
    .o(al_a1c88bcd));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*~(B)+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(B)+~(D)*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B)"),
    .INIT(32'h04378cbf))
    al_6f839cf3 (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_677d00f0[11]),
    .d(al_32c99495[11]),
    .e(al_42381c95[11]),
    .o(al_4a8487b2));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(~D*A))"),
    .INIT(16'h0cae))
    al_978656d6 (
    .a(al_f4b9a391),
    .b(al_e2aa4ae4),
    .c(al_a1c88bcd),
    .d(al_4a8487b2),
    .o(al_4197a0a2[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_3b570948 (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[12]),
    .o(al_a100d2c5[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hc3dff3dfcfdfffdf))
    al_22be5e53 (
    .a(al_a100d2c5[12]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .e(al_3cae1837[12]),
    .f(al_1cb63986[12]),
    .o(al_852e5bbe));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*~(B)+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(B)+~(D)*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B)"),
    .INIT(32'h04378cbf))
    al_18a823ab (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_677d00f0[12]),
    .d(al_32c99495[12]),
    .e(al_42381c95[12]),
    .o(al_ee5f9e50));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(~D*A))"),
    .INIT(16'h0cae))
    al_8234e90b (
    .a(al_f4b9a391),
    .b(al_e2aa4ae4),
    .c(al_852e5bbe),
    .d(al_ee5f9e50),
    .o(al_4197a0a2[12]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c047d0f4 (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[13]),
    .o(al_a100d2c5[13]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hc3dff3dfcfdfffdf))
    al_fcc38952 (
    .a(al_a100d2c5[13]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .e(al_3cae1837[13]),
    .f(al_1cb63986[13]),
    .o(al_1c6af38a));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*~(B)+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(B)+~(D)*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B)"),
    .INIT(32'h04378cbf))
    al_aa9fe077 (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_677d00f0[13]),
    .d(al_32c99495[13]),
    .e(al_42381c95[13]),
    .o(al_b3550f8b));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(~D*A))"),
    .INIT(16'h0cae))
    al_f350c8f3 (
    .a(al_f4b9a391),
    .b(al_e2aa4ae4),
    .c(al_1c6af38a),
    .d(al_b3550f8b),
    .o(al_4197a0a2[13]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f2a75e68 (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[14]),
    .o(al_a100d2c5[14]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hc3dff3dfcfdfffdf))
    al_6f2f506e (
    .a(al_a100d2c5[14]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .e(al_3cae1837[14]),
    .f(al_1cb63986[14]),
    .o(al_60adcd8c));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*~(B)+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(B)+~(D)*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B)"),
    .INIT(32'h04378cbf))
    al_fc694f5f (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_677d00f0[14]),
    .d(al_32c99495[14]),
    .e(al_42381c95[14]),
    .o(al_618a5a5f));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(~D*A))"),
    .INIT(16'h0cae))
    al_622816ba (
    .a(al_f4b9a391),
    .b(al_e2aa4ae4),
    .c(al_60adcd8c),
    .d(al_618a5a5f),
    .o(al_4197a0a2[14]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_44c46ea6 (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[15]),
    .o(al_a100d2c5[15]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hc3dff3dfcfdfffdf))
    al_e4238ee5 (
    .a(al_a100d2c5[15]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .e(al_3cae1837[15]),
    .f(al_1cb63986[15]),
    .o(al_1883a4da));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*~(B)+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(B)+~(D)*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B)"),
    .INIT(32'h04378cbf))
    al_1260f46e (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_677d00f0[15]),
    .d(al_32c99495[15]),
    .e(al_42381c95[15]),
    .o(al_f947ca8));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(~D*A))"),
    .INIT(16'h0cae))
    al_546d5029 (
    .a(al_f4b9a391),
    .b(al_e2aa4ae4),
    .c(al_1883a4da),
    .d(al_f947ca8),
    .o(al_4197a0a2[15]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_ed5691b1 (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[16]),
    .e(al_32c99495[16]),
    .f(al_42381c95[16]),
    .o(al_4197a0a2[16]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_5b15dc52 (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[17]),
    .e(al_32c99495[17]),
    .f(al_42381c95[17]),
    .o(al_4197a0a2[17]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_1f544b8 (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[18]),
    .e(al_32c99495[18]),
    .f(al_42381c95[18]),
    .o(al_4197a0a2[18]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_f1b27b9e (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[19]),
    .e(al_32c99495[19]),
    .f(al_42381c95[19]),
    .o(al_4197a0a2[19]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h236f))
    al_4441ef16 (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[7]),
    .c(al_871e6587[1]),
    .d(al_3cae1837[1]),
    .o(al_66a27b74));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~((E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*~((~D*~C))+~A*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)*~((~D*~C))+~(~A)*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)*(~D*~C)+~A*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)*(~D*~C))"),
    .INIT(64'haaa0aaa3aaacaaaf))
    al_81880382 (
    .a(al_66a27b74),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_eb5eeaf9[7]),
    .e(al_a3c2ad2a[1]),
    .f(al_44560df6[1]),
    .o(al_69ac11ac));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d4b2d82f (
    .a(al_eb5eeaf9[4]),
    .b(al_677d00f0[1]),
    .c(al_42381c95[1]),
    .o(al_52b0078[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfbf8cbc83b380b08))
    al_85c3bf4 (
    .a(al_52b0078[1]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[7]),
    .d(al_32c99495[1]),
    .e(al_3f753490[1]),
    .f(al_1cb63986[1]),
    .o(al_e340ee08[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .INIT(16'h44c0))
    al_5de6dfe1 (
    .a(al_69ac11ac),
    .b(al_e2aa4ae4),
    .c(al_e340ee08[1]),
    .d(al_eb5eeaf9[6]),
    .o(al_4197a0a2[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_57efa2e6 (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[20]),
    .e(al_32c99495[20]),
    .f(al_42381c95[20]),
    .o(al_4197a0a2[20]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_472197b (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[21]),
    .e(al_32c99495[21]),
    .f(al_42381c95[21]),
    .o(al_4197a0a2[21]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_d885e31b (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[22]),
    .e(al_32c99495[22]),
    .f(al_42381c95[22]),
    .o(al_4197a0a2[22]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_256fcbf7 (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[23]),
    .e(al_32c99495[23]),
    .f(al_42381c95[23]),
    .o(al_4197a0a2[23]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_2ad51b72 (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[24]),
    .e(al_32c99495[24]),
    .f(al_42381c95[24]),
    .o(al_4197a0a2[24]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_f30106ed (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[25]),
    .e(al_32c99495[25]),
    .f(al_42381c95[25]),
    .o(al_4197a0a2[25]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_9341608c (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[26]),
    .e(al_32c99495[26]),
    .f(al_42381c95[26]),
    .o(al_4197a0a2[26]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_8dc424f8 (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[27]),
    .e(al_32c99495[27]),
    .f(al_42381c95[27]),
    .o(al_4197a0a2[27]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_10203b04 (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[28]),
    .e(al_32c99495[28]),
    .f(al_42381c95[28]),
    .o(al_4197a0a2[28]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_716c7412 (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[29]),
    .e(al_32c99495[29]),
    .f(al_42381c95[29]),
    .o(al_4197a0a2[29]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_793de3ff (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[2]),
    .o(al_a100d2c5[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_673432e4 (
    .a(al_a100d2c5[2]),
    .b(al_eb5eeaf9[6]),
    .c(al_eb5eeaf9[7]),
    .d(al_32c99495[2]),
    .e(al_3f753490[2]),
    .f(al_3cae1837[2]),
    .o(al_36260f8d));
  AL_MAP_LUT6 #(
    .EQN("(~B*((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(F)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*F*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*F*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*F*C))"),
    .INIT(64'h3332313003020100))
    al_3b1aa32b (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[6]),
    .c(al_eb5eeaf9[7]),
    .d(al_677d00f0[2]),
    .e(al_42381c95[2]),
    .f(al_1cb63986[2]),
    .o(al_1d55dde3));
  AL_MAP_LUT4 #(
    .EQN("(A*(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D))"),
    .INIT(16'ha022))
    al_7432c9e2 (
    .a(al_e2aa4ae4),
    .b(al_36260f8d),
    .c(al_1d55dde3),
    .d(al_eb5eeaf9[5]),
    .o(al_4197a0a2[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_d4c51a3e (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[30]),
    .e(al_32c99495[30]),
    .f(al_42381c95[30]),
    .o(al_4197a0a2[30]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_293ebefa (
    .a(al_e2aa4ae4),
    .b(al_eb5eeaf9[6]),
    .c(al_eb5eeaf9[7]),
    .o(al_f4b9a391));
  AL_MAP_LUT6 #(
    .EQN("(A*(E*~((D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B))*~(C)+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*~(C)+~(E)*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C+E*(D*~(F)*~(B)+D*F*~(B)+~(D)*F*B+D*F*B)*C))"),
    .INIT(64'haa8aa0802a0a2000))
    al_71e85922 (
    .a(al_f4b9a391),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_677d00f0[31]),
    .e(al_32c99495[31]),
    .f(al_42381c95[31]),
    .o(al_4197a0a2[31]));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    al_2a560948 (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[7]),
    .c(al_a3c2ad2a[3]),
    .d(al_3cae1837[3]),
    .o(al_488ce459));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'he0efe3efecefefef))
    al_9f5ef007 (
    .a(al_488ce459),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .e(al_3f753490[3]),
    .f(al_1cb63986[3]),
    .o(al_2acb5425));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*~(B)+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(B)+~(D)*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B)"),
    .INIT(32'h04378cbf))
    al_28417d00 (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_677d00f0[3]),
    .d(al_32c99495[3]),
    .e(al_42381c95[3]),
    .o(al_8e73257f));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(~D*A))"),
    .INIT(16'h0cae))
    al_3bca93ca (
    .a(al_f4b9a391),
    .b(al_e2aa4ae4),
    .c(al_2acb5425),
    .d(al_8e73257f),
    .o(al_4197a0a2[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_57f9e609 (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[4]),
    .o(al_a100d2c5[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h04073437c4c7f4f7))
    al_e636bcc9 (
    .a(al_a100d2c5[4]),
    .b(al_eb5eeaf9[6]),
    .c(al_eb5eeaf9[7]),
    .d(al_32c99495[4]),
    .e(al_3f753490[4]),
    .f(al_3cae1837[4]),
    .o(al_5ecd0d98));
  AL_MAP_LUT6 #(
    .EQN("(~B*((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(F)*~(C)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*F*~(C)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*F*C+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*F*C))"),
    .INIT(64'h3332313003020100))
    al_bd99529d (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[6]),
    .c(al_eb5eeaf9[7]),
    .d(al_677d00f0[4]),
    .e(al_42381c95[4]),
    .f(al_1cb63986[4]),
    .o(al_b809a0d));
  AL_MAP_LUT4 #(
    .EQN("(A*(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D))"),
    .INIT(16'ha022))
    al_36b89aab (
    .a(al_e2aa4ae4),
    .b(al_5ecd0d98),
    .c(al_b809a0d),
    .d(al_eb5eeaf9[5]),
    .o(al_4197a0a2[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8cb504a9 (
    .a(al_eb5eeaf9[4]),
    .b(al_677d00f0[5]),
    .c(al_42381c95[5]),
    .o(al_52b0078[5]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfbf8cbc83b380b08))
    al_d246c0aa (
    .a(al_52b0078[5]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[7]),
    .d(al_32c99495[5]),
    .e(al_3f753490[5]),
    .f(al_1cb63986[5]),
    .o(al_e340ee08[5]));
  AL_MAP_LUT5 #(
    .EQN("(~B*((D*~A)*~(E)*~(C)+(D*~A)*E*~(C)+~((D*~A))*E*C+(D*~A)*E*C))"),
    .INIT(32'h31300100))
    al_f4c2372a (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[7]),
    .d(al_a3c2ad2a[5]),
    .e(al_3cae1837[5]),
    .o(al_9e3bc263[5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    al_f2d0fa8a (
    .a(al_e2aa4ae4),
    .b(al_e340ee08[5]),
    .c(al_9e3bc263[5]),
    .d(al_eb5eeaf9[6]),
    .o(al_4197a0a2[5]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_37dfb170 (
    .a(al_eb5eeaf9[0]),
    .b(al_eb5eeaf9[1]),
    .c(al_eb5eeaf9[2]),
    .d(al_eb5eeaf9[3]),
    .o(al_8b7519f2));
  AL_MAP_LUT5 #(
    .EQN("(B*(~A*~((~D*~C))*~(E)+~A*(~D*~C)*~(E)+~(~A)*(~D*~C)*E+~A*(~D*~C)*E))"),
    .INIT(32'h000c4444))
    al_4c09223 (
    .a(al_4db0ca34),
    .b(al_e2aa4ae4),
    .c(al_39575073),
    .d(al_eb5eeaf9[5]),
    .e(al_eb5eeaf9[6]),
    .o(al_4197a0a2[6]));
  AL_MAP_LUT5 #(
    .EQN("(A*(B*~(C)*~(D)*~(E)+~(B)*C*~(D)*~(E)+B*C*~(D)*~(E)+~(B)*~(C)*D*~(E)+B*~(C)*D*~(E)+~(B)*C*D*~(E)+B*C*D*~(E)+B*~(C)*~(D)*E+B*C*~(D)*E+~(B)*~(C)*D*E))"),
    .INIT(32'h0288aaa8))
    al_16ec2423 (
    .a(al_8b7519f2),
    .b(al_eb5eeaf9[4]),
    .c(al_eb5eeaf9[5]),
    .d(al_eb5eeaf9[6]),
    .e(al_eb5eeaf9[7]),
    .o(al_e2aa4ae4));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_ea84f218 (
    .a(al_3f753490[0]),
    .b(al_3f753490[1]),
    .c(al_3f753490[2]),
    .d(al_3f753490[3]),
    .e(al_3f753490[4]),
    .f(al_3f753490[5]),
    .o(al_46dd4bfb));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_5b2d8018 (
    .a(al_46dd4bfb),
    .b(al_3f753490[6]),
    .o(al_ec112ad9));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2d7862fc (
    .a(al_eb5eeaf9[4]),
    .b(al_677d00f0[6]),
    .c(al_42381c95[6]),
    .o(al_52b0078[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F)"),
    .INIT(64'h0530053ff530f53f))
    al_1835572f (
    .a(al_ec112ad9),
    .b(al_52b0078[6]),
    .c(al_eb5eeaf9[5]),
    .d(al_eb5eeaf9[7]),
    .e(al_32c99495[6]),
    .f(al_1cb63986[6]),
    .o(al_4db0ca34));
  AL_MAP_LUT4 #(
    .EQN("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .INIT(16'h23ef))
    al_cfb3a2f1 (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[7]),
    .c(al_a3c2ad2a[6]),
    .d(al_3cae1837[6]),
    .o(al_39575073));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d59557e (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[7]),
    .o(al_a100d2c5[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hc3dff3dfcfdfffdf))
    al_66455621 (
    .a(al_a100d2c5[7]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .e(al_3cae1837[7]),
    .f(al_1cb63986[7]),
    .o(al_f423313d));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*~(B)+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(B)+~(D)*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B)"),
    .INIT(32'h04378cbf))
    al_ad4d22f8 (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_677d00f0[7]),
    .d(al_32c99495[7]),
    .e(al_42381c95[7]),
    .o(al_ef0c62ea));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(~D*A))"),
    .INIT(16'h0cae))
    al_693d07ca (
    .a(al_f4b9a391),
    .b(al_e2aa4ae4),
    .c(al_f423313d),
    .d(al_ef0c62ea),
    .o(al_4197a0a2[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b70f9e23 (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[8]),
    .o(al_a100d2c5[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hc3dff3dfcfdfffdf))
    al_59bc8937 (
    .a(al_a100d2c5[8]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .e(al_3cae1837[8]),
    .f(al_1cb63986[8]),
    .o(al_56e2186e));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*~(B)+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(B)+~(D)*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B)"),
    .INIT(32'h04378cbf))
    al_c57996a (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_677d00f0[8]),
    .d(al_32c99495[8]),
    .e(al_42381c95[8]),
    .o(al_9e23e23c));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(~D*A))"),
    .INIT(16'h0cae))
    al_cfbf4ec1 (
    .a(al_f4b9a391),
    .b(al_e2aa4ae4),
    .c(al_56e2186e),
    .d(al_9e23e23c),
    .o(al_4197a0a2[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_8a445ab7 (
    .a(al_eb5eeaf9[4]),
    .b(al_a3c2ad2a[9]),
    .o(al_a100d2c5[9]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hc3dff3dfcfdfffdf))
    al_4fe2be21 (
    .a(al_a100d2c5[9]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .e(al_3cae1837[9]),
    .f(al_1cb63986[9]),
    .o(al_6cc2d7f5));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A))*~(B)+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*~(B)+~(D)*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B+D*(C*~(E)*~(A)+C*E*~(A)+~(C)*E*A+C*E*A)*B)"),
    .INIT(32'h04378cbf))
    al_aafac6e9 (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_677d00f0[9]),
    .d(al_32c99495[9]),
    .e(al_42381c95[9]),
    .o(al_71411c23));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(~D*A))"),
    .INIT(16'h0cae))
    al_90b3b0b3 (
    .a(al_f4b9a391),
    .b(al_e2aa4ae4),
    .c(al_6cc2d7f5),
    .d(al_71411c23),
    .o(al_4197a0a2[9]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_cf3eae0e (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[0]),
    .d(s_axi_wdata[0]),
    .e(al_42381c95[0]),
    .o(al_ae69e57d[0]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_54cc1f7c (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[10]),
    .d(s_axi_wdata[10]),
    .e(al_42381c95[10]),
    .o(al_ae69e57d[10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_c82b6db8 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[11]),
    .d(s_axi_wdata[11]),
    .e(al_42381c95[11]),
    .o(al_ae69e57d[11]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_474b95b6 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[12]),
    .d(s_axi_wdata[12]),
    .e(al_42381c95[12]),
    .o(al_ae69e57d[12]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_cc06f669 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[13]),
    .d(s_axi_wdata[13]),
    .e(al_42381c95[13]),
    .o(al_ae69e57d[13]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_932e93a2 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[14]),
    .d(s_axi_wdata[14]),
    .e(al_42381c95[14]),
    .o(al_ae69e57d[14]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_5fc9f079 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[15]),
    .d(s_axi_wdata[15]),
    .e(al_42381c95[15]),
    .o(al_ae69e57d[15]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_6e2b046f (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[16]),
    .d(s_axi_wdata[16]),
    .e(al_42381c95[16]),
    .o(al_ae69e57d[16]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_161734f9 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[17]),
    .d(s_axi_wdata[17]),
    .e(al_42381c95[17]),
    .o(al_ae69e57d[17]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_de103e2b (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[18]),
    .d(s_axi_wdata[18]),
    .e(al_42381c95[18]),
    .o(al_ae69e57d[18]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_993a03ff (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[19]),
    .d(s_axi_wdata[19]),
    .e(al_42381c95[19]),
    .o(al_ae69e57d[19]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_5baaa7e4 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[1]),
    .d(s_axi_wdata[1]),
    .e(al_42381c95[1]),
    .o(al_ae69e57d[1]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_70d0a6 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[20]),
    .d(s_axi_wdata[20]),
    .e(al_42381c95[20]),
    .o(al_ae69e57d[20]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_69a738bf (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[21]),
    .d(s_axi_wdata[21]),
    .e(al_42381c95[21]),
    .o(al_ae69e57d[21]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_f2443a0b (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[22]),
    .d(s_axi_wdata[22]),
    .e(al_42381c95[22]),
    .o(al_ae69e57d[22]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_c5d16ebb (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[23]),
    .d(s_axi_wdata[23]),
    .e(al_42381c95[23]),
    .o(al_ae69e57d[23]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_81f0670f (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[24]),
    .d(s_axi_wdata[24]),
    .e(al_42381c95[24]),
    .o(al_ae69e57d[24]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_3e8ad80b (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[25]),
    .d(s_axi_wdata[25]),
    .e(al_42381c95[25]),
    .o(al_ae69e57d[25]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_6b13715f (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[26]),
    .d(s_axi_wdata[26]),
    .e(al_42381c95[26]),
    .o(al_ae69e57d[26]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_2f2f0867 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[27]),
    .d(s_axi_wdata[27]),
    .e(al_42381c95[27]),
    .o(al_ae69e57d[27]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_e5b2e9bb (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[28]),
    .d(s_axi_wdata[28]),
    .e(al_42381c95[28]),
    .o(al_ae69e57d[28]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_c4fc65ba (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[29]),
    .d(s_axi_wdata[29]),
    .e(al_42381c95[29]),
    .o(al_ae69e57d[29]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_29846a32 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[2]),
    .d(s_axi_wdata[2]),
    .e(al_42381c95[2]),
    .o(al_ae69e57d[2]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_8ae1da87 (
    .a(al_9daabc69),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_b93f6564));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_eedecab6 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[30]),
    .d(s_axi_wdata[30]),
    .e(al_42381c95[30]),
    .o(al_ae69e57d[30]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_8824e8f8 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[31]),
    .d(s_axi_wdata[31]),
    .e(al_42381c95[31]),
    .o(al_ae69e57d[31]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_fc7f3471 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[3]),
    .d(s_axi_wdata[3]),
    .e(al_42381c95[3]),
    .o(al_ae69e57d[3]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_dbd52179 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[4]),
    .d(s_axi_wdata[4]),
    .e(al_42381c95[4]),
    .o(al_ae69e57d[4]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_6ff332a3 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[5]),
    .d(s_axi_wdata[5]),
    .e(al_42381c95[5]),
    .o(al_ae69e57d[5]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_41476af2 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[6]),
    .d(s_axi_wdata[6]),
    .e(al_42381c95[6]),
    .o(al_ae69e57d[6]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_9975b0fb (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[7]),
    .d(s_axi_wdata[7]),
    .e(al_42381c95[7]),
    .o(al_ae69e57d[7]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_c00ced96 (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[8]),
    .d(s_axi_wdata[8]),
    .e(al_42381c95[8]),
    .o(al_ae69e57d[8]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_fae64a7f (
    .a(al_b93f6564),
    .b(al_655c284a),
    .c(pause_source_addr[9]),
    .d(s_axi_wdata[9]),
    .e(al_42381c95[9]),
    .o(al_ae69e57d[9]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_fa9e39a9 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[32]),
    .d(s_axi_wdata[0]),
    .e(al_a3c2ad2a[0]),
    .o(al_1062ede0[0]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_60e6df29 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[42]),
    .d(s_axi_wdata[10]),
    .e(al_a3c2ad2a[10]),
    .o(al_1062ede0[10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_82fe9a92 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[43]),
    .d(s_axi_wdata[11]),
    .e(al_a3c2ad2a[11]),
    .o(al_1062ede0[11]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_7446f4e6 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[44]),
    .d(s_axi_wdata[12]),
    .e(al_a3c2ad2a[12]),
    .o(al_1062ede0[12]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_83780304 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[45]),
    .d(s_axi_wdata[13]),
    .e(al_a3c2ad2a[13]),
    .o(al_1062ede0[13]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_d60efa04 (
    .a(al_16296d60),
    .b(al_677d00f0[0]),
    .o(al_655c284a));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*~B*A)"),
    .INIT(32'h00000200))
    al_5c9341de (
    .a(al_9daabc69),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_e1f066de));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_439664c0 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[46]),
    .d(s_axi_wdata[14]),
    .e(al_a3c2ad2a[14]),
    .o(al_1062ede0[14]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_f533bad5 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[47]),
    .d(s_axi_wdata[15]),
    .e(al_a3c2ad2a[15]),
    .o(al_1062ede0[15]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_49093e53 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[33]),
    .d(s_axi_wdata[1]),
    .e(al_a3c2ad2a[1]),
    .o(al_1062ede0[1]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_e7b3a7d9 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[34]),
    .d(s_axi_wdata[2]),
    .e(al_a3c2ad2a[2]),
    .o(al_1062ede0[2]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_f0a82cb (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[35]),
    .d(s_axi_wdata[3]),
    .e(al_a3c2ad2a[3]),
    .o(al_1062ede0[3]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_818c60a8 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[36]),
    .d(s_axi_wdata[4]),
    .e(al_a3c2ad2a[4]),
    .o(al_1062ede0[4]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_8bde4ede (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[37]),
    .d(s_axi_wdata[5]),
    .e(al_a3c2ad2a[5]),
    .o(al_1062ede0[5]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_83532cbf (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[38]),
    .d(s_axi_wdata[6]),
    .e(al_a3c2ad2a[6]),
    .o(al_1062ede0[6]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_63ba75bf (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[39]),
    .d(s_axi_wdata[7]),
    .e(al_a3c2ad2a[7]),
    .o(al_1062ede0[7]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_f9db84c4 (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[40]),
    .d(s_axi_wdata[8]),
    .e(al_a3c2ad2a[8]),
    .o(al_1062ede0[8]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_28ecf66a (
    .a(al_e1f066de),
    .b(al_655c284a),
    .c(pause_source_addr[41]),
    .d(s_axi_wdata[9]),
    .e(al_a3c2ad2a[9]),
    .o(al_1062ede0[9]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_cd1ee769 (
    .a(al_16296d60),
    .b(al_32c99495[0]),
    .o(al_7fda1410));
  AL_DFF_0 al_2955d836 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9d802914),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0936433));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(A)*~((F*E*~C))+D*A*~((F*E*~C))+~(D)*A*(F*E*~C)+D*A*(F*E*~C)))"),
    .INIT(64'h3202330033003300))
    al_3e7b3189 (
    .a(al_ec112ad9),
    .b(al_16296d60),
    .c(al_86bf0006),
    .d(al_c0936433),
    .e(al_8bef06bd),
    .f(al_a15918b4),
    .o(al_9d802914));
  AL_DFF_0 al_db1d817c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_86bf0006),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_8bef06bd));
  AL_DFF_0 al_62bfd959 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(mdio_in),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_27629aac));
  AL_DFF_0 al_d90a5adc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_27629aac),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_3560f04f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F)"),
    .INIT(64'h555533330f0f00ff))
    al_d07aec3c (
    .a(al_3cae1837[8]),
    .b(al_3cae1837[9]),
    .c(al_3cae1837[10]),
    .d(al_3cae1837[11]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_6a277bd4));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F)"),
    .INIT(64'h555533330f0f00ff))
    al_ddf89d40 (
    .a(al_3cae1837[0]),
    .b(al_3cae1837[1]),
    .c(al_3cae1837[2]),
    .d(al_3cae1837[3]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_f1c0fe91));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00ccccf0f0aaaa))
    al_e433c003 (
    .a(al_27f7f6ec),
    .b(al_afd5fd5d),
    .c(al_6a277bd4),
    .d(al_f1c0fe91),
    .e(al_71b90bfa[2]),
    .f(al_71b90bfa[3]),
    .o(al_18128b53));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h33330f0f00ff5555))
    al_5549992d (
    .a(al_7de51101[3]),
    .b(al_7de51101[10]),
    .c(al_7de51101[11]),
    .d(al_7de51101[12]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_12c9315c));
  AL_MAP_LUT6 #(
    .EQN("~(~(~(B)*~(C)*D*~(E)+B*~(C)*D*~(E)+~(B)*C*D*~(E)+B*C*D*~(E)+~(B)*C*~(D)*E+B*C*~(D)*E+B*~(C)*D*E+B*C*D*E)*~(A)*~(F)+~(~(B)*~(C)*D*~(E)+B*~(C)*D*~(E)+~(B)*C*D*~(E)+B*C*D*~(E)+~(B)*C*~(D)*E+B*C*~(D)*E+B*~(C)*D*E+B*C*D*E)*A*~(F)+~(~(~(B)*~(C)*D*~(E)+B*~(C)*D*~(E)+~(B)*C*D*~(E)+B*C*D*~(E)+~(B)*C*~(D)*E+B*C*~(D)*E+B*~(C)*D*E+B*C*D*E))*A*F+~(~(B)*~(C)*D*~(E)+B*~(C)*D*~(E)+~(B)*C*D*~(E)+B*C*D*~(E)+~(B)*C*~(D)*E+B*C*~(D)*E+B*~(C)*D*E+B*C*D*E)*A*F)"),
    .INIT(64'h55555555ccf0ff00))
    al_71c294c0 (
    .a(al_12c9315c),
    .b(al_7de51101[1]),
    .c(al_7de51101[2]),
    .d(al_71b90bfa[0]),
    .e(al_71b90bfa[1]),
    .f(al_71b90bfa[3]),
    .o(al_54829ae8));
  AL_DFF_0 al_142a2a0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_830d7e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mdio_out));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F)"),
    .INIT(64'h555533330f0f00ff))
    al_15de4d59 (
    .a(al_7de51101[4]),
    .b(al_7de51101[5]),
    .c(al_7de51101[6]),
    .d(al_7de51101[7]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_7360a7c0));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((~(B)*C*~(D)*~(E)+B*C*~(D)*~(E)+B*~(C)*D*~(E)+B*C*D*~(E)+~(B)*~(C)*~(D)*E+B*~(C)*~(D)*E+~(B)*C*~(D)*E+B*C*~(D)*E))*~(F)+~A*(~(B)*C*~(D)*~(E)+B*C*~(D)*~(E)+B*~(C)*D*~(E)+B*C*D*~(E)+~(B)*~(C)*~(D)*E+B*~(C)*~(D)*E+~(B)*C*~(D)*E+B*C*~(D)*E)*~(F)+~(~A)*(~(B)*C*~(D)*~(E)+B*C*~(D)*~(E)+B*~(C)*D*~(E)+B*C*D*~(E)+~(B)*~(C)*~(D)*E+B*~(C)*~(D)*E+~(B)*C*~(D)*E+B*C*~(D)*E)*F+~A*(~(B)*C*~(D)*~(E)+B*C*~(D)*~(E)+B*~(C)*D*~(E)+B*C*D*~(E)+~(B)*~(C)*~(D)*E+B*~(C)*~(D)*E+~(B)*C*~(D)*E+B*C*~(D)*E)*F)"),
    .INIT(64'h00ffccf055555555))
    al_8ca23264 (
    .a(al_7360a7c0),
    .b(al_7de51101[8]),
    .c(al_7de51101[9]),
    .d(al_71b90bfa[0]),
    .e(al_71b90bfa[1]),
    .f(al_71b90bfa[3]),
    .o(al_5cbbf9cd));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(A)*~(E)+~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*~(E)+~(~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*A*E+~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*E)"),
    .INIT(32'haaaa0f33))
    al_1b123f43 (
    .a(al_18128b53),
    .b(al_54829ae8),
    .c(al_5cbbf9cd),
    .d(al_71b90bfa[2]),
    .e(al_71b90bfa[4]),
    .o(al_2d86aa6e));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(~E*~((F*A))*~((D*~C))+~E*(F*A)*~((D*~C))+~(~E)*(F*A)*(D*~C)+~E*(F*A)*(D*~C)))"),
    .INIT(64'h3133010033330300))
    al_6bc96c7c (
    .a(al_2d86aa6e),
    .b(al_16296d60),
    .c(al_86bf0006),
    .d(al_8bef06bd),
    .e(mdio_out),
    .f(al_71b90bfa[5]),
    .o(al_830d7e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F)"),
    .INIT(64'h555533330f0f00ff))
    al_7997239f (
    .a(al_3cae1837[12]),
    .b(al_3cae1837[13]),
    .c(al_3cae1837[14]),
    .d(al_3cae1837[15]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_27f7f6ec));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F)"),
    .INIT(64'h555533330f0f00ff))
    al_d11f65b3 (
    .a(al_3cae1837[4]),
    .b(al_3cae1837[5]),
    .c(al_3cae1837[6]),
    .d(al_3cae1837[7]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_afd5fd5d));
  AL_DFF_1 al_3960090e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_63df2227),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mdio_oen));
  AL_MAP_LUT6 #(
    .EQN("(F*A*~(~E*~(D*C*B)))"),
    .INIT(64'haaaa800000000000))
    al_d38bc0b (
    .a(al_7de51101[2]),
    .b(al_71b90bfa[1]),
    .c(al_71b90bfa[2]),
    .d(al_71b90bfa[3]),
    .e(al_71b90bfa[4]),
    .f(al_71b90bfa[5]),
    .o(al_12b617e9));
  AL_MAP_LUT6 #(
    .EQN("~(~B*(~E*~((~F*~A))*~((D*~C))+~E*(~F*~A)*~((D*~C))+~(~E)*(~F*~A)*(D*~C)+~E*(~F*~A)*(D*~C)))"),
    .INIT(64'hffffcfccfeffcecc))
    al_17589ec0 (
    .a(al_12b617e9),
    .b(al_16296d60),
    .c(al_86bf0006),
    .d(al_8bef06bd),
    .e(mdio_oen),
    .f(al_a15918b4),
    .o(al_63df2227));
  AL_DFF_1 al_ffed6b0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_aecc1a53),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a15918b4));
  AL_MAP_LUT6 #(
    .EQN("~(~C*(~(A)*~(B)*~((E*D))*~(F)+A*~(B)*~((E*D))*~(F)+~(A)*B*~((E*D))*~(F)+~(A)*~(B)*(E*D)*~(F)+A*~(B)*(E*D)*~(F)+~(A)*B*(E*D)*~(F)+~(A)*B*(E*D)*F))"),
    .INIT(64'hfbfffffff8f8f8f8))
    al_58409d35 (
    .a(al_77c268d4),
    .b(al_ae3e538d),
    .c(al_16296d60),
    .d(al_1ff3d4e5),
    .e(al_c0936433),
    .f(al_a15918b4),
    .o(al_aecc1a53));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_340a0cbe (
    .a(al_ae3e538d),
    .b(al_71b90bfa[2]),
    .c(al_71b90bfa[3]),
    .d(al_71b90bfa[4]),
    .e(al_71b90bfa[5]),
    .o(al_5d42041c));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((F*~E*A))+D*C*~((F*~E*A))+~(D)*C*(F*~E*A)+D*C*(F*~E*A)))"),
    .INIT(64'h3300312033003300))
    al_c33b3ced (
    .a(al_5d42041c),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[1]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_6492ae8));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((~F*E*A))+D*C*~((~F*E*A))+~(D)*C*(~F*E*A)+D*C*(~F*E*A)))"),
    .INIT(64'h3300330031203300))
    al_3935c4b7 (
    .a(al_5d42041c),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[2]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_9e9040d4));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((~F*~E*A))+D*C*~((~F*~E*A))+~(D)*C*(~F*~E*A)+D*C*(~F*~E*A)))"),
    .INIT(64'h3300330033003120))
    al_c7118da4 (
    .a(al_5d42041c),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[3]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_f44ba8da));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*A)"),
    .INIT(32'h20000000))
    al_c4897809 (
    .a(al_ae3e538d),
    .b(al_71b90bfa[2]),
    .c(al_71b90bfa[3]),
    .d(al_71b90bfa[4]),
    .e(al_71b90bfa[5]),
    .o(al_f78634c8));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((F*E*A))+D*C*~((F*E*A))+~(D)*C*(F*E*A)+D*C*(F*E*A)))"),
    .INIT(64'h3120330033003300))
    al_1309f9a5 (
    .a(al_f78634c8),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[4]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_adf2eefc));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((F*~E*A))+D*C*~((F*~E*A))+~(D)*C*(F*~E*A)+D*C*(F*~E*A)))"),
    .INIT(64'h3300312033003300))
    al_360897e0 (
    .a(al_f78634c8),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[5]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_944f1baf));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((~F*E*A))+D*C*~((~F*E*A))+~(D)*C*(~F*E*A)+D*C*(~F*E*A)))"),
    .INIT(64'h3300330031203300))
    al_a6d3b535 (
    .a(al_f78634c8),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[6]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_ee5a9fb));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((~F*~E*A))+D*C*~((~F*~E*A))+~(D)*C*(~F*~E*A)+D*C*(~F*~E*A)))"),
    .INIT(64'h3300330033003120))
    al_30bcfead (
    .a(al_f78634c8),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[7]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_15e31402));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*B*A)"),
    .INIT(32'h08000000))
    al_a2600967 (
    .a(al_ae3e538d),
    .b(al_71b90bfa[2]),
    .c(al_71b90bfa[3]),
    .d(al_71b90bfa[4]),
    .e(al_71b90bfa[5]),
    .o(al_33d9db52));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((F*E*A))+D*C*~((F*E*A))+~(D)*C*(F*E*A)+D*C*(F*E*A)))"),
    .INIT(64'h3120330033003300))
    al_9013b123 (
    .a(al_33d9db52),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[8]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_955255ce));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((F*~E*A))+D*C*~((F*~E*A))+~(D)*C*(F*~E*A)+D*C*(F*~E*A)))"),
    .INIT(64'h3300312033003300))
    al_1fb62a49 (
    .a(al_33d9db52),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[9]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_61af39ad));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((~F*E*A))+D*C*~((~F*E*A))+~(D)*C*(~F*E*A)+D*C*(~F*E*A)))"),
    .INIT(64'h3300330031203300))
    al_7e52faee (
    .a(al_33d9db52),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[10]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_20afe6c0));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((~F*~E*A))+D*C*~((~F*~E*A))+~(D)*C*(~F*~E*A)+D*C*(~F*~E*A)))"),
    .INIT(64'h3300330033003120))
    al_61cc7d82 (
    .a(al_33d9db52),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[11]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_138eaec3));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*A)"),
    .INIT(32'h02000000))
    al_fbd594ff (
    .a(al_ae3e538d),
    .b(al_71b90bfa[2]),
    .c(al_71b90bfa[3]),
    .d(al_71b90bfa[4]),
    .e(al_71b90bfa[5]),
    .o(al_6b647f54));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((F*E*A))+D*C*~((F*E*A))+~(D)*C*(F*E*A)+D*C*(F*E*A)))"),
    .INIT(64'h3120330033003300))
    al_f9ce3fb (
    .a(al_6b647f54),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[12]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_72045a1c));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((F*~E*A))+D*C*~((F*~E*A))+~(D)*C*(F*~E*A)+D*C*(F*~E*A)))"),
    .INIT(64'h3300312033003300))
    al_1eba92d7 (
    .a(al_6b647f54),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[13]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_ee917930));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((~F*E*A))+D*C*~((~F*E*A))+~(D)*C*(~F*E*A)+D*C*(~F*E*A)))"),
    .INIT(64'h3300330031203300))
    al_28b957b4 (
    .a(al_6b647f54),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[14]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_88c12a03));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((~F*~E*A))+D*C*~((~F*~E*A))+~(D)*C*(~F*~E*A)+D*C*(~F*~E*A)))"),
    .INIT(64'h3300330033003120))
    al_aef55aa9 (
    .a(al_6b647f54),
    .b(al_16296d60),
    .c(al_3560f04f),
    .d(al_1cb63986[15]),
    .e(al_71b90bfa[0]),
    .f(al_71b90bfa[1]),
    .o(al_ddac5e8d));
  AL_DFF_0 al_42eabff (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_46fb2129),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[0]));
  AL_DFF_0 al_2be91d7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6492ae8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[1]));
  AL_DFF_0 al_ed37bfb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9e9040d4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[2]));
  AL_DFF_0 al_4c5fd1b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_f44ba8da),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[3]));
  AL_DFF_0 al_cca4168d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_adf2eefc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[4]));
  AL_DFF_0 al_d202e609 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_944f1baf),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[5]));
  AL_DFF_0 al_e7748593 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ee5a9fb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[6]));
  AL_DFF_0 al_8501cec4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_15e31402),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[7]));
  AL_DFF_0 al_9765c304 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_955255ce),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[8]));
  AL_DFF_0 al_abd07723 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_61af39ad),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[9]));
  AL_DFF_0 al_b23a06c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_20afe6c0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[10]));
  AL_DFF_0 al_a56f6eae (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_138eaec3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[11]));
  AL_DFF_0 al_4b4c65ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_72045a1c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[12]));
  AL_DFF_0 al_bfa465e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ee917930),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[13]));
  AL_DFF_0 al_31eb251e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_88c12a03),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[14]));
  AL_DFF_0 al_d6cae29c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddac5e8d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1cb63986[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_6ec51051 (
    .a(al_7f161bf2),
    .b(al_71b90bfa[4]),
    .c(al_71b90bfa[5]),
    .o(al_77c268d4));
  AL_MAP_LUT5 #(
    .EQN("(~C*(E*~(D)*~((B*A))+E*D*~((B*A))+~(E)*D*(B*A)+E*D*(B*A)))"),
    .INIT(32'h0f070800))
    al_8ecdfbfd (
    .a(al_77c268d4),
    .b(al_ae3e538d),
    .c(al_16296d60),
    .d(al_3560f04f),
    .e(al_1cb63986[0]),
    .o(al_46fb2129));
  AL_DFF_0 al_78bee461 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_fabf91f7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71b90bfa[2]));
  AL_DFF_0 al_90d8b017 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_2169fa2d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71b90bfa[3]));
  AL_DFF_0 al_ea23f275 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_a698f8f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71b90bfa[4]));
  AL_DFF_0 al_faf3c9d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_14067aef),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71b90bfa[5]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_35c72738 (
    .a(al_71b90bfa[0]),
    .b(al_71b90bfa[1]),
    .c(al_71b90bfa[2]),
    .d(al_71b90bfa[3]),
    .o(al_7f161bf2));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_c7ba226f (
    .a(al_86bf0006),
    .b(al_8bef06bd),
    .o(al_ae3e538d));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(C)*~(D)+~(A)*~(C)*D+~(A)*C*D))"),
    .INIT(16'h1102))
    al_c9312861 (
    .a(al_ae3e538d),
    .b(al_16296d60),
    .c(al_a15918b4),
    .d(al_71b90bfa[0]),
    .o(al_c3ba6eaa));
  AL_MAP_LUT5 #(
    .EQN("(~B*(A*~(C)*D*~(E)+~(A)*~(C)*~(D)*E+A*~(C)*~(D)*E+~(A)*C*~(D)*E+~(A)*~(C)*D*E+~(A)*C*D*E))"),
    .INIT(32'h11130200))
    al_b40d86f0 (
    .a(al_ae3e538d),
    .b(al_16296d60),
    .c(al_a15918b4),
    .d(al_71b90bfa[0]),
    .e(al_71b90bfa[1]),
    .o(al_338b9100));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*(E*D)*~(F)+~(A)*~(C)*~((E*D))*F+A*~(C)*~((E*D))*F+~(A)*C*~((E*D))*F+~(A)*~(C)*(E*D)*F+~(A)*C*(E*D)*F))"),
    .INIT(64'h1113131302000000))
    al_55886208 (
    .a(al_ae3e538d),
    .b(al_16296d60),
    .c(al_a15918b4),
    .d(al_71b90bfa[0]),
    .e(al_71b90bfa[1]),
    .f(al_71b90bfa[2]),
    .o(al_fabf91f7));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_c06eb13b (
    .a(al_71b90bfa[0]),
    .b(al_71b90bfa[1]),
    .c(al_71b90bfa[2]),
    .o(al_4f925611));
  AL_MAP_LUT5 #(
    .EQN("(~C*(A*B*~(D)*~(E)+~(A)*~(B)*~(D)*E+A*~(B)*~(D)*E+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*~(B)*D*E))"),
    .INIT(32'h03070008))
    al_ba6108b2 (
    .a(al_4f925611),
    .b(al_ae3e538d),
    .c(al_16296d60),
    .d(al_a15918b4),
    .e(al_71b90bfa[3]),
    .o(al_2169fa2d));
  AL_MAP_LUT5 #(
    .EQN("(~C*(A*B*~(D)*~(E)+~(A)*~(B)*~(D)*E+A*~(B)*~(D)*E+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*~(B)*D*E))"),
    .INIT(32'h03070008))
    al_d6aa77e3 (
    .a(al_7f161bf2),
    .b(al_ae3e538d),
    .c(al_16296d60),
    .d(al_a15918b4),
    .e(al_71b90bfa[4]),
    .o(al_a698f8f));
  AL_MAP_LUT6 #(
    .EQN("(~C*(B*~(D)*(E*A)*~(F)+~(B)*~(D)*~((E*A))*F+B*~(D)*~((E*A))*F+~(B)*D*~((E*A))*F+~(B)*~(D)*(E*A)*F+~(B)*D*(E*A)*F))"),
    .INIT(64'h0307030f00080000))
    al_754a331f (
    .a(al_7f161bf2),
    .b(al_ae3e538d),
    .c(al_16296d60),
    .d(al_a15918b4),
    .e(al_71b90bfa[4]),
    .f(al_71b90bfa[5]),
    .o(al_14067aef));
  AL_DFF_0 al_a665fc8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_c3ba6eaa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71b90bfa[0]));
  AL_DFF_0 al_872ed2a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_338b9100),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_71b90bfa[1]));
  AL_DFF_0 al_1e33afd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_77c268d4),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_60f51d47));
  AL_DFF_0 al_157dc1ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_60f51d47),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_9439ddc));
  AL_DFF_X al_68728a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d7a47bf6),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_18642257));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_76974295 (
    .a(al_cc7e79c9),
    .b(al_e1057698),
    .o(al_41d2ce29));
  AL_DFF_X al_fb5eb836 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_41d2ce29),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_a37dea2d));
  AL_DFF_X al_11fef992 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b3220547),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_39c05299));
  AL_MAP_LUT5 #(
    .EQN("(~E*(D*~(C)*~((B*A))+D*C*~((B*A))+~(D)*C*(B*A)+D*C*(B*A)))"),
    .INIT(32'h0000f780))
    al_668f7120 (
    .a(al_6f75ef0e),
    .b(rx_clk_en),
    .c(al_677d00f0[4]),
    .d(al_39c05299),
    .e(al_fea77e50),
    .o(al_b3220547));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_2897c6e6 (
    .a(al_583c216b[0]),
    .b(al_583c216b[2]),
    .c(al_583c216b[4]),
    .d(al_583c216b[6]),
    .e(al_583c216b[7]),
    .o(al_8f689368));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(~F*~E*~D*~C*A))"),
    .INIT(64'h3333333333333331))
    al_cbc7cfd5 (
    .a(al_8f689368),
    .b(al_dd43c64f),
    .c(al_7a7628f9),
    .d(al_583c216b[1]),
    .e(al_583c216b[3]),
    .f(al_583c216b[5]),
    .o(al_d6baa558));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b16cbcfa (
    .a(al_d6baa558),
    .b(al_d83e61fb),
    .o(al_1bdd94f8));
  AL_DFF_X al_2ced7a17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1bdd94f8),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_dd43c64f));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_7098fd (
    .a(al_4c1d19df),
    .b(al_cc7e79c9),
    .c(al_7ac96e46),
    .o(al_9a2dcc24));
  AL_DFF_X al_fe01963a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9a2dcc24),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_c2520419));
  AL_DFF_0 al_8698ddf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_bf03de15),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81b839ee[0]));
  AL_DFF_0 al_9b07cfcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_81b839ee[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81b839ee[1]));
  AL_DFF_0 al_ba6b8769 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_81b839ee[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81b839ee[2]));
  AL_DFF_0 al_50c50519 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_81b839ee[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81b839ee[3]));
  AL_DFF_0 al_89a1da02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_81b839ee[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81b839ee[4]));
  AL_DFF_0 al_70cb5cd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_81b839ee[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81b839ee[5]));
  AL_DFF_0 al_83b892c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_932a07c7),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_469f2a04[0]));
  AL_DFF_0 al_11074846 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_469f2a04[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_469f2a04[1]));
  AL_DFF_0 al_e2cd01e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_469f2a04[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_469f2a04[2]));
  AL_DFF_0 al_78b60c81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7a7628f9),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff43a01c[0]));
  AL_DFF_0 al_2c7f4ac1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ff43a01c[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff43a01c[1]));
  AL_DFF_0 al_ae4de999 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ff43a01c[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff43a01c[2]));
  AL_DFF_0 al_47eb96f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ff43a01c[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff43a01c[3]));
  AL_DFF_X al_1b32f23f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_677d00f0[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_4c9b2533));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_efedf4c0 (
    .a(al_1d03242c[2]),
    .b(al_1d03242c[3]),
    .c(al_1d03242c[4]),
    .d(al_1d03242c[5]),
    .e(al_1d03242c[6]),
    .f(al_1d03242c[7]),
    .o(al_7710deab));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*A)"),
    .INIT(32'h20000000))
    al_27bcb9b6 (
    .a(al_7710deab),
    .b(al_62730356),
    .c(al_ebdfe328),
    .d(al_1d03242c[0]),
    .e(al_1d03242c[1]),
    .o(al_4696ac48));
  AL_DFF_X al_c7807a50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4696ac48),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_c5450b82));
  AL_DFF_X al_4dea5c5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9809ce8b),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_6e672ebc));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_dfedc68b (
    .a(rx_clk_en),
    .b(al_4c9b2533),
    .o(al_e890f462));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_6758468e (
    .a(al_124e348a),
    .b(al_1a0f7d2b[0]),
    .c(al_fdc321a5),
    .o(al_e57de54[0]));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*A))"),
    .INIT(8'h6c))
    al_b1fef4e6 (
    .a(al_b70fe470),
    .b(al_53a2c384[2]),
    .c(al_fdc321a5),
    .o(al_e57de54[10]));
  AL_MAP_LUT6 #(
    .EQN("(D@(F*(E@C@B@A)))"),
    .INIT(64'h96696996ff00ff00))
    al_d64d245c (
    .a(al_5107a44a),
    .b(al_d9299255),
    .c(al_1a0f7d2b[7]),
    .d(al_53a2c384[3]),
    .e(al_53a2c384[24]),
    .f(al_fdc321a5),
    .o(al_e57de54[11]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_422b407b (
    .a(al_d671f8ef),
    .b(al_f00de1fc),
    .o(al_b605ded6));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*(C@B@A)))"),
    .INIT(32'h6996ff00))
    al_5e3ebd4f (
    .a(al_b605ded6),
    .b(al_124e348a),
    .c(al_d9299255),
    .d(al_53a2c384[4]),
    .e(al_fdc321a5),
    .o(al_e57de54[12]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_682b737d (
    .a(al_1a0f7d2b[5]),
    .b(al_53a2c384[26]),
    .o(al_f00de1fc));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_390d3611 (
    .a(al_1a0f7d2b[1]),
    .b(al_1a0f7d2b[2]),
    .c(al_53a2c384[29]),
    .d(al_53a2c384[30]),
    .o(al_4409fb45));
  AL_MAP_LUT6 #(
    .EQN("(E@(F*(D@C@B@A)))"),
    .INIT(64'h96696996ffff0000))
    al_2399812a (
    .a(al_e34977fd),
    .b(al_4409fb45),
    .c(al_a3a88d3f),
    .d(al_f00de1fc),
    .e(al_53a2c384[5]),
    .f(al_fdc321a5),
    .o(al_e57de54[13]));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    al_d630062c (
    .a(al_a3a88d3f),
    .b(al_1a0f7d2b[3]),
    .c(al_53a2c384[28]),
    .o(al_5107a44a));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*~(C@B@A)))"),
    .INIT(32'h9669ff00))
    al_90425614 (
    .a(al_5107a44a),
    .b(al_5f1c4763[0]),
    .c(al_f00de1fc),
    .d(al_53a2c384[6]),
    .e(al_fdc321a5),
    .o(al_e57de54[14]));
  AL_MAP_LUT6 #(
    .EQN("(D@(F*(E@C@B@A)))"),
    .INIT(64'h96696996ff00ff00))
    al_58b24a1c (
    .a(al_d671f8ef),
    .b(al_a3a88d3f),
    .c(al_1a0f7d2b[0]),
    .d(al_53a2c384[7]),
    .e(al_53a2c384[31]),
    .f(al_fdc321a5),
    .o(al_e57de54[15]));
  AL_MAP_LUT5 #(
    .EQN("(C@(E*~(D@B@A)))"),
    .INIT(32'h9669f0f0))
    al_b3591822 (
    .a(al_d671f8ef),
    .b(al_1a0f7d2b[7]),
    .c(al_53a2c384[8]),
    .d(al_53a2c384[24]),
    .e(al_fdc321a5),
    .o(al_e57de54[16]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*~(B@A)))"),
    .INIT(16'h69f0))
    al_ad0b214a (
    .a(al_4409fb45),
    .b(al_d9299255),
    .c(al_53a2c384[9]),
    .d(al_fdc321a5),
    .o(al_e57de54[17]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*~(B@A)))"),
    .INIT(16'h69f0))
    al_b2329455 (
    .a(al_5f1c4763[0]),
    .b(al_f00de1fc),
    .c(al_53a2c384[10]),
    .d(al_fdc321a5),
    .o(al_e57de54[18]));
  AL_MAP_LUT5 #(
    .EQN("(C@(E*(D@B@A)))"),
    .INIT(32'h6996f0f0))
    al_20571e80 (
    .a(al_a3a88d3f),
    .b(al_1a0f7d2b[0]),
    .c(al_53a2c384[11]),
    .d(al_53a2c384[31]),
    .e(al_fdc321a5),
    .o(al_e57de54[19]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_7dab301d (
    .a(al_c611b356),
    .b(al_1a0f7d2b[1]),
    .c(al_fdc321a5),
    .o(al_e57de54[1]));
  AL_MAP_LUT4 #(
    .EQN("(B@(D*~(C@A)))"),
    .INIT(16'h69cc))
    al_3d9f42b0 (
    .a(al_1a0f7d2b[3]),
    .b(al_53a2c384[12]),
    .c(al_53a2c384[28]),
    .d(al_fdc321a5),
    .o(al_e57de54[20]));
  AL_MAP_LUT4 #(
    .EQN("(B@(D*~(C@A)))"),
    .INIT(16'h69cc))
    al_27ed006 (
    .a(al_1a0f7d2b[2]),
    .b(al_53a2c384[13]),
    .c(al_53a2c384[29]),
    .d(al_fdc321a5),
    .o(al_e57de54[21]));
  AL_MAP_LUT4 #(
    .EQN("(B@(D*~(C@A)))"),
    .INIT(16'h69cc))
    al_5ffe0d66 (
    .a(al_1a0f7d2b[7]),
    .b(al_53a2c384[14]),
    .c(al_53a2c384[24]),
    .d(al_fdc321a5),
    .o(al_e57de54[22]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*~(B@A)))"),
    .INIT(16'h69f0))
    al_1af6cd98 (
    .a(al_124e348a),
    .b(al_d9299255),
    .c(al_53a2c384[15]),
    .d(al_fdc321a5),
    .o(al_e57de54[23]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*~(B@A)))"),
    .INIT(16'h69f0))
    al_214efce5 (
    .a(al_e34977fd),
    .b(al_f00de1fc),
    .c(al_53a2c384[16]),
    .d(al_fdc321a5),
    .o(al_e57de54[24]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*(B@A)))"),
    .INIT(16'h96f0))
    al_23aac1e7 (
    .a(al_a3a88d3f),
    .b(al_f00de1fc),
    .c(al_53a2c384[17]),
    .d(al_fdc321a5),
    .o(al_e57de54[25]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*(B@A)))"),
    .INIT(16'h96f0))
    al_5c71c91b (
    .a(al_5107a44a),
    .b(al_124e348a),
    .c(al_53a2c384[18]),
    .d(al_fdc321a5),
    .o(al_e57de54[26]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*(B@A)))"),
    .INIT(16'h96f0))
    al_c98496f6 (
    .a(al_e34977fd),
    .b(al_d671f8ef),
    .c(al_53a2c384[19]),
    .d(al_fdc321a5),
    .o(al_e57de54[27]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*~(B@A)))"),
    .INIT(16'h69f0))
    al_699dbcf6 (
    .a(al_4409fb45),
    .b(al_f00de1fc),
    .c(al_53a2c384[20]),
    .d(al_fdc321a5),
    .o(al_e57de54[28]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*~(B@A)))"),
    .INIT(16'h69f0))
    al_9accec7 (
    .a(al_5f1c4763[0]),
    .b(al_a3a88d3f),
    .c(al_53a2c384[21]),
    .d(al_fdc321a5),
    .o(al_e57de54[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~((B@A))*~(D)+C*(B@A)*~(D)+~(C)*(B@A)*D+C*(B@A)*D)"),
    .INIT(16'h66f0))
    al_6cafef58 (
    .a(al_c611b356),
    .b(al_f00de1fc),
    .c(al_1a0f7d2b[2]),
    .d(al_fdc321a5),
    .o(al_e57de54[2]));
  AL_MAP_LUT6 #(
    .EQN("(C@(F*(E@D@B@A)))"),
    .INIT(64'h96696996f0f0f0f0))
    al_cb8bae5b (
    .a(al_1a0f7d2b[0]),
    .b(al_1a0f7d2b[3]),
    .c(al_53a2c384[22]),
    .d(al_53a2c384[28]),
    .e(al_53a2c384[31]),
    .f(al_fdc321a5),
    .o(al_e57de54[30]));
  AL_MAP_LUT4 #(
    .EQN("(B@(D*~(C@A)))"),
    .INIT(16'h69cc))
    al_ddf35a20 (
    .a(al_1a0f7d2b[2]),
    .b(al_53a2c384[23]),
    .c(al_53a2c384[29]),
    .d(al_fdc321a5),
    .o(al_e57de54[31]));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~((C@B@A))*~(E)+~D*(C@B@A)*~(E)+~(~D)*(C@B@A)*E+~D*(C@B@A)*E)"),
    .INIT(32'h6969ff00))
    al_ab376a8e (
    .a(al_e34977fd),
    .b(al_a3a88d3f),
    .c(al_f00de1fc),
    .d(al_1a0f7d2b[3]),
    .e(al_fdc321a5),
    .o(al_e57de54[3]));
  AL_MAP_LUT5 #(
    .EQN("(D*~((C@B@A))*~(E)+D*(C@B@A)*~(E)+~(D)*(C@B@A)*E+D*(C@B@A)*E)"),
    .INIT(32'h9696ff00))
    al_eab5e43e (
    .a(al_5107a44a),
    .b(al_124e348a),
    .c(al_f00de1fc),
    .d(al_1a0f7d2b[4]),
    .e(al_fdc321a5),
    .o(al_e57de54[4]));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_c847a468 (
    .a(al_1a0f7d2b[1]),
    .b(al_1a0f7d2b[7]),
    .c(al_53a2c384[24]),
    .d(al_53a2c384[30]),
    .o(al_124e348a));
  AL_MAP_LUT5 #(
    .EQN("(D*~((C@B@A))*~(E)+D*(C@B@A)*~(E)+~(D)*(C@B@A)*E+D*(C@B@A)*E)"),
    .INIT(32'h9696ff00))
    al_e9a24adf (
    .a(al_c611b356),
    .b(al_d671f8ef),
    .c(al_a3a88d3f),
    .d(al_1a0f7d2b[5]),
    .e(al_fdc321a5),
    .o(al_e57de54[5]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_5619eee6 (
    .a(al_1a0f7d2b[4]),
    .b(al_53a2c384[27]),
    .o(al_a3a88d3f));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_35e7ee1c (
    .a(al_1a0f7d2b[6]),
    .b(al_53a2c384[25]),
    .o(al_d9299255));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_60546d75 (
    .a(al_1a0f7d2b[2]),
    .b(al_1a0f7d2b[3]),
    .c(al_53a2c384[28]),
    .d(al_53a2c384[29]),
    .o(al_d671f8ef));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    al_dcc5a0f (
    .a(al_d9299255),
    .b(al_1a0f7d2b[0]),
    .c(al_53a2c384[31]),
    .o(al_e34977fd));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_ae2d8e78 (
    .a(al_e34977fd),
    .b(al_124e348a),
    .o(al_c611b356));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_ee2a4b2a (
    .a(al_1a0f7d2b[0]),
    .b(al_1a0f7d2b[1]),
    .c(al_53a2c384[30]),
    .d(al_53a2c384[31]),
    .o(al_5f1c4763[0]));
  AL_MAP_LUT5 #(
    .EQN("(C@(E*~(D@B@A)))"),
    .INIT(32'h9669f0f0))
    al_28c500d5 (
    .a(al_b605ded6),
    .b(al_5f1c4763[0]),
    .c(al_1a0f7d2b[6]),
    .d(al_53a2c384[25]),
    .e(al_fdc321a5),
    .o(al_e57de54[6]));
  AL_MAP_LUT6 #(
    .EQN("(F@E@D@C@B@A)"),
    .INIT(64'h6996966996696996))
    al_a1e328cb (
    .a(al_a3a88d3f),
    .b(al_f00de1fc),
    .c(al_1a0f7d2b[2]),
    .d(al_1a0f7d2b[7]),
    .e(al_53a2c384[24]),
    .f(al_53a2c384[29]),
    .o(al_b70fe470));
  AL_MAP_LUT5 #(
    .EQN("(C*~((D@B@A))*~(E)+C*(D@B@A)*~(E)+~(C)*(D@B@A)*E+C*(D@B@A)*E)"),
    .INIT(32'h9966f0f0))
    al_b5a60831 (
    .a(al_b70fe470),
    .b(al_1a0f7d2b[0]),
    .c(al_1a0f7d2b[7]),
    .d(al_53a2c384[31]),
    .e(al_fdc321a5),
    .o(al_e57de54[7]));
  AL_MAP_LUT6 #(
    .EQN("(D@(F*(E@C@B@A)))"),
    .INIT(64'h96696996ff00ff00))
    al_1c95e7d6 (
    .a(al_5107a44a),
    .b(al_d9299255),
    .c(al_1a0f7d2b[7]),
    .d(al_53a2c384[0]),
    .e(al_53a2c384[24]),
    .f(al_fdc321a5),
    .o(al_e57de54[8]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*(B@A)))"),
    .INIT(16'h96f0))
    al_f23aa978 (
    .a(al_b605ded6),
    .b(al_d9299255),
    .c(al_53a2c384[1]),
    .d(al_fdc321a5),
    .o(al_e57de54[9]));
  AL_DFF_X al_3362c12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[8]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[8]));
  AL_DFF_X al_ebc2c67b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[9]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[9]));
  AL_DFF_X al_3e70e048 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[10]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[10]));
  AL_DFF_X al_24671ab7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[11]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[11]));
  AL_DFF_X al_270484bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[12]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[12]));
  AL_DFF_X al_f76e6f06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[13]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[13]));
  AL_DFF_X al_e87aef22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[14]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[14]));
  AL_DFF_X al_c943323 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[15]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[15]));
  AL_DFF_X al_1693b7df (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[16]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[16]));
  AL_DFF_X al_4b101b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[17]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[17]));
  AL_DFF_X al_36d539e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[0]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[0]));
  AL_DFF_X al_db06c75f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[18]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[18]));
  AL_DFF_X al_a77d0094 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[19]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[19]));
  AL_DFF_X al_c3f345c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[20]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[20]));
  AL_DFF_X al_b833f575 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[21]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[21]));
  AL_DFF_X al_882784b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[22]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[22]));
  AL_DFF_X al_9781d129 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[23]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[23]));
  AL_DFF_X al_70366825 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[24]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[24]));
  AL_DFF_X al_1d606cf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[25]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[25]));
  AL_DFF_X al_f868a692 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[26]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[26]));
  AL_DFF_X al_97b486c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[27]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[27]));
  AL_DFF_X al_2bfe74eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[1]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[1]));
  AL_DFF_X al_8fdc0b43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[28]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[28]));
  AL_DFF_X al_eb3f2b49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[29]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[29]));
  AL_DFF_X al_6a84056f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[30]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[30]));
  AL_DFF_X al_925d72e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[31]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[31]));
  AL_DFF_X al_88d87aad (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[2]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[2]));
  AL_DFF_X al_a0c808f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[3]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[3]));
  AL_DFF_X al_f527cce3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[4]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[4]));
  AL_DFF_X al_1af1fb14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[5]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[5]));
  AL_DFF_X al_2cc8a9ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[6]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[6]));
  AL_DFF_X al_4303127 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e57de54[7]),
    .en(al_e890f462),
    .sr(al_6f75ef0e),
    .ss(1'b0),
    .q(al_53a2c384[7]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*~A))"),
    .INIT(16'h00fe))
    al_723960b6 (
    .a(al_e78cfe9),
    .b(al_aceaab6b),
    .c(al_d7a47bf6),
    .d(al_5d14a06f),
    .o(al_8b0ea091));
  AL_DFF_X al_a95cc281 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8b0ea091),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_d7a47bf6));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~E*~D*~C*~A))"),
    .INIT(32'hccccccc8))
    al_e820597 (
    .a(al_2eea7a5a),
    .b(al_ce4327dc),
    .c(al_36b29f2),
    .d(al_decf41ac),
    .e(al_81378cfb),
    .o(al_f0d27177));
  AL_DFF_X al_5f227e09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0d27177),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e1057698));
  AL_MAP_LUT6 #(
    .EQN("(~(D@C)*~(E@B)*~(F@A))"),
    .INIT(64'h8008200240041001))
    al_134b2b7d (
    .a(al_1a0f7d2b[2]),
    .b(al_1a0f7d2b[3]),
    .c(al_1a0f7d2b[7]),
    .d(al_53a2c384[24]),
    .e(al_53a2c384[28]),
    .f(al_53a2c384[29]),
    .o(al_bbbfb344));
  AL_MAP_LUT5 #(
    .EQN("(~C*~B*A*~(E@D))"),
    .INIT(32'h02000002))
    al_234f0d45 (
    .a(al_bbbfb344),
    .b(al_a3a88d3f),
    .c(al_f00de1fc),
    .d(al_1a0f7d2b[1]),
    .e(al_53a2c384[30]),
    .o(al_66f2b6b8));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~B*A*~(D@C)))"),
    .INIT(32'hdffd0000))
    al_d516f47d (
    .a(al_66f2b6b8),
    .b(al_d9299255),
    .c(al_1a0f7d2b[0]),
    .d(al_53a2c384[31]),
    .e(al_a409c88e),
    .o(al_46839cba));
  AL_DFF_X al_111c3472 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_46839cba),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_13cf5eba));
  AL_DFF_X al_275f5e8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2eea7a5a),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e5a67968));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*B)))"),
    .INIT(16'h00ea))
    al_d07129e (
    .a(al_f3170c9),
    .b(al_45a6c91),
    .c(al_e2dc2eea),
    .d(al_5d14a06f),
    .o(al_2270269f));
  AL_DFF_X al_d0aaa631 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2270269f),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f3170c9));
  AL_DFF_X al_ca8acd6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8fc9814c),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_179ef786));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    al_82eaae1d (
    .a(al_2eea7a5a),
    .b(al_7ffbbf6e),
    .c(al_7c1aee64),
    .d(al_db678397),
    .o(al_1fad8912));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(D*~B)))"),
    .INIT(16'h0705))
    al_2dddab26 (
    .a(al_1fad8912),
    .b(al_c5450b82),
    .c(al_5d14a06f),
    .d(al_8fc9814c),
    .o(al_ba6d5331));
  AL_DFF_X al_d0698bd1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ba6d5331),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_df30c316));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D*B)))"),
    .INIT(16'hbafa))
    al_6d6a3d8d (
    .a(al_88bee87),
    .b(al_179ef786),
    .c(al_38e61a96),
    .d(al_db678397),
    .o(al_43d0de98));
  AL_DFF_X al_20149c83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_43d0de98),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_38e61a96));
  AL_MAP_LUT6 #(
    .EQN("(~(D*~C)*~(~(E*~B)*~(F*~A)))"),
    .INIT(64'h7077505530330000))
    al_82c18e8a (
    .a(al_74c05d28),
    .b(al_6c6d3d88),
    .c(al_f3170c9),
    .d(al_45a6c91),
    .e(al_1ce99d34),
    .f(al_8c3b9f16),
    .o(al_12dfe9dc));
  AL_MAP_LUT6 #(
    .EQN("(F*~(~A*~(~E*~D*~C*~B)))"),
    .INIT(64'haaaaaaab00000000))
    al_f1da7e4c (
    .a(al_12dfe9dc),
    .b(al_74c05d28),
    .c(al_dacf8588),
    .d(al_8c3b9f16),
    .e(al_31cc16da),
    .f(al_4d5dd241),
    .o(al_75def4ef));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~C*~A*~(D*~B)))"),
    .INIT(32'h0000fbfa))
    al_234ec4b6 (
    .a(al_75def4ef),
    .b(al_f3170c9),
    .c(al_36b29f2),
    .d(al_a409c88e),
    .e(al_5d14a06f),
    .o(al_d4a11187));
  AL_DFF_X al_15489660 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d4a11187),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36b29f2));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_83c97354 (
    .a(al_13cf5eba),
    .b(al_df30c316),
    .o(al_2eea7a5a));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_539a1203 (
    .a(al_134f4cf5),
    .b(al_5d14a06f),
    .o(al_ce4327dc));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*~A)"),
    .INIT(32'h00000004))
    al_5061c8f6 (
    .a(al_2eea7a5a),
    .b(al_ce4327dc),
    .c(al_36b29f2),
    .d(al_decf41ac),
    .e(al_81378cfb),
    .o(al_aa9f8872));
  AL_DFF_X al_4606a227 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aa9f8872),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_d6bd6336));
  AL_DFF_X al_9a011a05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_153d6f9e),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_44348d99));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    al_57bc28d6 (
    .a(al_6f75ef0e),
    .b(al_134f4cf5),
    .c(al_5d14a06f),
    .o(al_21b2c715));
  AL_DFF_X al_d8df8251 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_21b2c715),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_134f4cf5));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_6619cda (
    .a(al_36b29f2),
    .b(al_31cc16da),
    .o(al_49b1129));
  AL_DFF_X al_e8deaaa9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_49b1129),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_b95885c7));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*D*~C*B*~A)"),
    .INIT(64'h0000040000000000))
    al_14779365 (
    .a(al_1e120105[0]),
    .b(al_1e120105[1]),
    .c(al_1e120105[4]),
    .d(al_1e120105[5]),
    .e(al_1e120105[9]),
    .f(al_1e120105[10]),
    .o(al_c4d37b2));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*~C*~(~B*A))"),
    .INIT(64'h0d00000000000000))
    al_eb90b438 (
    .a(al_3ccf053a),
    .b(al_1e120105[2]),
    .c(al_1e120105[3]),
    .d(al_1e120105[6]),
    .e(al_1e120105[7]),
    .f(al_1e120105[8]),
    .o(al_1dcf5c5b));
  AL_MAP_LUT6 #(
    .EQN("(~E*~C*~(~D*~(~F*B*A)))"),
    .INIT(64'h00000f0000000f08))
    al_8b1013c0 (
    .a(al_c4d37b2),
    .b(al_1dcf5c5b),
    .c(al_225d06ad),
    .d(al_decf41ac),
    .e(al_5d14a06f),
    .f(al_8fc9814c),
    .o(al_d49fbba9));
  AL_DFF_X al_8930e15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d49fbba9),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_decf41ac));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*~C*B*~A)"),
    .INIT(64'h0000000000000400))
    al_dbb46788 (
    .a(al_1e120105[0]),
    .b(al_1e120105[1]),
    .c(al_1e120105[4]),
    .d(al_1e120105[5]),
    .e(al_1e120105[6]),
    .f(al_1e120105[7]),
    .o(al_2ac16c9f));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_a0d23627 (
    .a(al_2ac16c9f),
    .b(al_1e120105[2]),
    .c(al_1e120105[3]),
    .o(al_7c20ee3b));
  AL_DFF_X al_d086285e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7c20ee3b),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_45a6c91));
  AL_DFF_X al_92e98474 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_decf41ac),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f5080327));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C@B))"),
    .INIT(8'hbe))
    al_711f6eff (
    .a(al_88bee87),
    .b(al_e9f83d6e),
    .c(al_e023302[0]),
    .o(al_5c2983f8[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(C*B)))"),
    .INIT(16'h1540))
    al_64d72aa1 (
    .a(al_88bee87),
    .b(al_e9f83d6e),
    .c(al_e023302[0]),
    .d(al_e023302[1]),
    .o(al_5c2983f8[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(E@(D*C*B)))"),
    .INIT(32'h15554000))
    al_f1257879 (
    .a(al_88bee87),
    .b(al_e9f83d6e),
    .c(al_e023302[0]),
    .d(al_e023302[1]),
    .e(al_e023302[2]),
    .o(al_5c2983f8[2]));
  AL_MAP_LUT6 #(
    .EQN("(~A*(F@(E*D*C*B)))"),
    .INIT(64'h1555555540000000))
    al_dea5d1a (
    .a(al_88bee87),
    .b(al_e9f83d6e),
    .c(al_e023302[0]),
    .d(al_e023302[1]),
    .e(al_e023302[2]),
    .f(al_e023302[3]),
    .o(al_5c2983f8[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_e06eb7dc (
    .a(al_88bee87),
    .b(al_9613edfd),
    .c(al_e023302[4]),
    .o(al_5c2983f8[4]));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_7e851e2 (
    .a(al_e9f83d6e),
    .b(al_e023302[0]),
    .c(al_e023302[1]),
    .d(al_e023302[2]),
    .e(al_e023302[3]),
    .o(al_9613edfd));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(C*B)))"),
    .INIT(16'h1540))
    al_5125f000 (
    .a(al_88bee87),
    .b(al_9613edfd),
    .c(al_e023302[4]),
    .d(al_e023302[5]),
    .o(al_5c2983f8[5]));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_3284e339 (
    .a(al_88bee87),
    .b(al_32ab2441),
    .c(al_e023302[6]),
    .o(al_5c2983f8[6]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(C*B)))"),
    .INIT(16'h1540))
    al_bf707232 (
    .a(al_88bee87),
    .b(al_32ab2441),
    .c(al_e023302[6]),
    .d(al_e023302[7]),
    .o(al_5c2983f8[7]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(E@(D*C*B)))"),
    .INIT(32'h15554000))
    al_b881b7b6 (
    .a(al_88bee87),
    .b(al_32ab2441),
    .c(al_e023302[6]),
    .d(al_e023302[7]),
    .e(al_e023302[8]),
    .o(al_5c2983f8[8]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_d71ac33a (
    .a(al_6b3de12e),
    .b(al_4f800f89),
    .c(al_db678397),
    .d(al_5b221454),
    .o(al_153d6f9e));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~F*~(E*D*C*B)))"),
    .INIT(64'h5555555540000000))
    al_b40224b (
    .a(al_88bee87),
    .b(al_32ab2441),
    .c(al_e023302[6]),
    .d(al_e023302[7]),
    .e(al_e023302[8]),
    .f(al_e023302[9]),
    .o(al_5c2983f8[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_65c3b0c4 (
    .a(al_153d6f9e),
    .b(al_44348d99),
    .o(al_88bee87));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e2ffc55b (
    .a(al_f02638e3),
    .b(al_e023302[6]),
    .c(al_e023302[9]),
    .o(al_c57a154));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(~F*~D*A*~(E*~C)))"),
    .INIT(64'h3333333333133311))
    al_50b48117 (
    .a(al_6b3de12e),
    .b(al_c57a154),
    .c(al_38e61a96),
    .d(al_4f800f89),
    .e(al_db678397),
    .f(al_5b221454),
    .o(al_e9f83d6e));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_cffd2c1 (
    .a(al_e023302[0]),
    .b(al_e023302[1]),
    .c(al_e023302[2]),
    .d(al_e023302[3]),
    .e(al_e023302[4]),
    .f(al_e023302[5]),
    .o(al_b610aa54));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_e60048e0 (
    .a(al_e9f83d6e),
    .b(al_b610aa54),
    .o(al_32ab2441));
  AL_MAP_LUT6 #(
    .EQN("(C*~(F*B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)))"),
    .INIT(64'h30b070f0f0f0f0f0))
    al_a20e764e (
    .a(al_f02638e3),
    .b(al_179ef786),
    .c(al_81378cfb),
    .d(al_7b9b882d[6]),
    .e(al_7b9b882d[9]),
    .f(al_db678397),
    .o(al_3f4108ac));
  AL_MAP_LUT6 #(
    .EQN("((B*~(~F*E*C))*~(D)*~(A)+(B*~(~F*E*C))*D*~(A)+~((B*~(~F*E*C)))*D*A+(B*~(~F*E*C))*D*A)"),
    .INIT(64'hee44ee44ae04ee44))
    al_f5212c26 (
    .a(al_88bee87),
    .b(al_3f4108ac),
    .c(al_c57a154),
    .d(al_9cabf6c6),
    .e(al_38e61a96),
    .f(al_db678397),
    .o(al_31415f80));
  AL_DFF_X al_6d711410 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_31415f80),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_81378cfb));
  AL_DFF_X al_5c2ce9a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ce4327dc),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_60b3be17));
  AL_DFF_X al_6292cdc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e023302[9]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7b9b882d[9]));
  AL_DFF_X al_d2e4889a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e023302[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7b9b882d[6]));
  AL_DFF_X al_db907b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5c2983f8[8]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e023302[8]));
  AL_DFF_X al_6396f757 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5c2983f8[9]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e023302[9]));
  AL_DFF_X al_b187fccd (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5c2983f8[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_e023302[0]));
  AL_DFF_X al_c5be1287 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5c2983f8[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e023302[1]));
  AL_DFF_X al_12a2d855 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5c2983f8[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e023302[2]));
  AL_DFF_X al_ebc890da (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5c2983f8[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e023302[3]));
  AL_DFF_X al_9a80eda3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5c2983f8[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e023302[4]));
  AL_DFF_X al_fbe8db0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5c2983f8[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e023302[5]));
  AL_DFF_X al_d1cec66e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5c2983f8[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e023302[6]));
  AL_DFF_X al_a9acd973 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5c2983f8[7]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e023302[7]));
  AL_MAP_LUT6 #(
    .EQN("(D*~C*~B*~A*~(~F*~E))"),
    .INIT(64'h0100010001000000))
    al_70d4dc42 (
    .a(al_1a0f7d2b[0]),
    .b(al_1a0f7d2b[1]),
    .c(al_1a0f7d2b[2]),
    .d(al_1a0f7d2b[3]),
    .e(al_484c4f9e),
    .f(al_3aba2254),
    .o(al_3e9eebf5));
  AL_MAP_LUT5 #(
    .EQN("((~E*C)*~((B*A))*~(D)+(~E*C)*(B*A)*~(D)+~((~E*C))*(B*A)*D+(~E*C)*(B*A)*D)"),
    .INIT(32'h880088f0))
    al_72b8800a (
    .a(al_3e9eebf5),
    .b(al_162f415f),
    .c(al_1e582b4d),
    .d(al_a468a88f),
    .e(al_5d14a06f),
    .o(al_9c659f6));
  AL_DFF_X al_65521864 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9c659f6),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e582b4d));
  AL_DFF_X al_ab8b5bce (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1e582b4d),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_384019b7));
  AL_DFF_X al_3037666e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_384019b7),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_b2deb19c));
  AL_MAP_LUT6 #(
    .EQN("(F*E*~D*~C*~B*A)"),
    .INIT(64'h0002000000000000))
    al_d9cc7726 (
    .a(al_162f415f),
    .b(al_1a0f7d2b[0]),
    .c(al_1a0f7d2b[1]),
    .d(al_1a0f7d2b[2]),
    .e(al_1a0f7d2b[3]),
    .f(al_a468a88f),
    .o(al_5c7d4b11));
  AL_MAP_LUT5 #(
    .EQN("((C*~B)*~(A)*~((E*D))+(C*~B)*A*~((E*D))+~((C*~B))*A*(E*D)+(C*~B)*A*(E*D))"),
    .INIT(32'haa303030))
    al_84ef66e9 (
    .a(al_5c7d4b11),
    .b(al_6f75ef0e),
    .c(al_abdbe49),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_b3d5e449));
  AL_DFF_X al_3728fc7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b3d5e449),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_abdbe49));
  AL_DFF_X al_73e40dac (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_abdbe49),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1ce99d34));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_63ebed3c (
    .a(al_4c3c2401),
    .b(al_1a0f7d2b[0]),
    .c(al_1a0f7d2b[1]),
    .d(al_1a0f7d2b[2]),
    .e(al_1a0f7d2b[3]),
    .o(al_ae1bb7ab));
  AL_DFF_X al_b28d1e1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ae1bb7ab),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_a468a88f));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(~D*~C*B))"),
    .INIT(16'haaae))
    al_a5ab3752 (
    .a(al_6f75ef0e),
    .b(al_fdc321a5),
    .c(al_4d5dd241),
    .d(al_5d14a06f),
    .o(al_bc9d849e));
  AL_DFF_X al_78b4cfa2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_bc9d849e),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_fdc321a5));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B@A))"),
    .INIT(8'h09))
    al_f5455958 (
    .a(al_6b3de12e),
    .b(al_1e120105[0]),
    .c(al_5d14a06f),
    .o(al_ea827a0c[0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_973e8509 (
    .a(al_a409c88e),
    .b(al_e2dc2eea),
    .c(al_8fc9814c),
    .d(al_fd106601),
    .o(al_6b3de12e));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_6df29789 (
    .a(al_6b3de12e),
    .b(al_1e120105[0]),
    .c(al_1e120105[1]),
    .o(al_30e55692));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_1a353e5b (
    .a(al_30e55692),
    .b(al_1e120105[2]),
    .c(al_1e120105[3]),
    .d(al_1e120105[4]),
    .e(al_1e120105[5]),
    .f(al_1e120105[6]),
    .o(al_efa05a0c));
  AL_MAP_LUT6 #(
    .EQN("(~F*(E@(D*C*B*A)))"),
    .INIT(64'h000000007fff8000))
    al_278b2cc2 (
    .a(al_efa05a0c),
    .b(al_1e120105[7]),
    .c(al_1e120105[8]),
    .d(al_1e120105[9]),
    .e(al_1e120105[10]),
    .f(al_5d14a06f),
    .o(al_ea827a0c[10]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C@(B*~A)))"),
    .INIT(16'h00b4))
    al_e1d3ff5 (
    .a(al_6b3de12e),
    .b(al_1e120105[0]),
    .c(al_1e120105[1]),
    .d(al_5d14a06f),
    .o(al_ea827a0c[1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*(B@A))"),
    .INIT(8'h06))
    al_c4d4b0b8 (
    .a(al_30e55692),
    .b(al_1e120105[2]),
    .c(al_5d14a06f),
    .o(al_ea827a0c[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C@(B*A)))"),
    .INIT(16'h0078))
    al_9f73368 (
    .a(al_30e55692),
    .b(al_1e120105[2]),
    .c(al_1e120105[3]),
    .d(al_5d14a06f),
    .o(al_ea827a0c[3]));
  AL_MAP_LUT5 #(
    .EQN("(~E*(D@(C*B*A)))"),
    .INIT(32'h00007f80))
    al_f8f23a93 (
    .a(al_30e55692),
    .b(al_1e120105[2]),
    .c(al_1e120105[3]),
    .d(al_1e120105[4]),
    .e(al_5d14a06f),
    .o(al_ea827a0c[4]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(E@(D*C*B*A)))"),
    .INIT(64'h000000007fff8000))
    al_b7de5f1f (
    .a(al_30e55692),
    .b(al_1e120105[2]),
    .c(al_1e120105[3]),
    .d(al_1e120105[4]),
    .e(al_1e120105[5]),
    .f(al_5d14a06f),
    .o(al_ea827a0c[5]));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_e423c186 (
    .a(al_30e55692),
    .b(al_1e120105[2]),
    .c(al_1e120105[3]),
    .d(al_1e120105[4]),
    .e(al_1e120105[5]),
    .f(al_1e120105[6]),
    .o(al_4f3b20c[6]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_335cebda (
    .a(al_4f3b20c[6]),
    .b(al_5d14a06f),
    .o(al_ea827a0c[6]));
  AL_MAP_LUT3 #(
    .EQN("(~C*(B@A))"),
    .INIT(8'h06))
    al_8de7657d (
    .a(al_efa05a0c),
    .b(al_1e120105[7]),
    .c(al_5d14a06f),
    .o(al_ea827a0c[7]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C@(B*A)))"),
    .INIT(16'h0078))
    al_7c4f8488 (
    .a(al_efa05a0c),
    .b(al_1e120105[7]),
    .c(al_1e120105[8]),
    .d(al_5d14a06f),
    .o(al_ea827a0c[8]));
  AL_MAP_LUT5 #(
    .EQN("(~E*(D@(C*B*A)))"),
    .INIT(32'h00007f80))
    al_37720fbf (
    .a(al_efa05a0c),
    .b(al_1e120105[7]),
    .c(al_1e120105[8]),
    .d(al_1e120105[9]),
    .e(al_5d14a06f),
    .o(al_ea827a0c[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_98449462 (
    .a(al_cb67e17c),
    .b(al_db678397),
    .o(al_6f75ef0e));
  AL_MAP_LUT5 #(
    .EQN("(~E*~C*~(~D*B*~A))"),
    .INIT(32'h00000f0b))
    al_580581e3 (
    .a(al_74c05d28),
    .b(al_dacf8588),
    .c(al_f9e26d2b),
    .d(al_31cc16da),
    .e(al_5d14a06f),
    .o(al_8a98fa0e));
  AL_MAP_LUT6 #(
    .EQN("~(~B*~(~D*C*A*~(F*E)))"),
    .INIT(64'hccccccecccecccec))
    al_8e7ee3e5 (
    .a(al_8a98fa0e),
    .b(al_6f75ef0e),
    .c(al_42c40cf0),
    .d(al_16c52309),
    .e(al_e2dc2eea),
    .f(al_4d5dd241),
    .o(al_a095939));
  AL_DFF_X al_626b1f49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_a095939),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_42c40cf0));
  AL_MAP_LUT6 #(
    .EQN("((~F*~E*~D*B)*~(C)*~(A)+(~F*~E*~D*B)*C*~(A)+~((~F*~E*~D*B))*C*A+(~F*~E*~D*B)*C*A)"),
    .INIT(64'ha0a0a0a0a0a0a0e4))
    al_f0fadfad (
    .a(al_39c05299),
    .b(al_42c40cf0),
    .c(al_9a3d38d8),
    .d(al_f9e26d2b),
    .e(al_5d14a06f),
    .f(al_8fc9814c),
    .o(al_df322506));
  AL_DFF_X al_2ac2992d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_df322506),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7ac96e46));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(~B*~A))"),
    .INIT(16'h0eee))
    al_5ffc390d (
    .a(al_6f75ef0e),
    .b(al_9a3d38d8),
    .c(al_a409c88e),
    .d(al_2c3ff84c),
    .o(al_ac4196c0));
  AL_DFF_X al_de79d749 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ac4196c0),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_9a3d38d8));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_1ac1b7ea (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[0]),
    .c(al_b9d3b2c1[0]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_179f9221 (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[10]),
    .c(al_b9d3b2c1[10]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[10]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_6a505a8 (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[11]),
    .c(al_b9d3b2c1[11]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[11]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_6dc6485d (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[12]),
    .c(al_b9d3b2c1[12]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[12]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_d4e71279 (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[13]),
    .c(al_b9d3b2c1[13]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[13]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    al_3163f8c7 (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[14]),
    .c(al_b9d3b2c1[14]),
    .o(al_9e843f7[14]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_e0e5acdc (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[1]),
    .c(al_b9d3b2c1[1]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[1]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_8fb134a4 (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[2]),
    .c(al_b9d3b2c1[2]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[2]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_3296d6ad (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[3]),
    .c(al_b9d3b2c1[3]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[3]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_92b1d17f (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[4]),
    .c(al_b9d3b2c1[4]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[4]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_81aa917c (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[5]),
    .c(al_b9d3b2c1[5]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[5]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_86a226b1 (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[6]),
    .c(al_b9d3b2c1[6]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[6]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_ab945a6a (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[7]),
    .c(al_b9d3b2c1[7]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[7]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_fbf85ba6 (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[8]),
    .c(al_b9d3b2c1[8]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[8]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_5269d206 (
    .a(al_6f75ef0e),
    .b(al_66bdfa10[9]),
    .c(al_b9d3b2c1[9]),
    .d(al_b9d3b2c1[14]),
    .o(al_9e843f7[9]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_421eee56 (
    .a(al_1e120105[1]),
    .b(al_1e120105[2]),
    .c(al_1e120105[3]),
    .d(al_2814a16d[1]),
    .e(al_2814a16d[2]),
    .f(al_2814a16d[3]),
    .o(al_13154bf6));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_6106ebcd (
    .a(al_b242277f),
    .b(al_5d14a06f),
    .o(al_509509ae));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_97db9118 (
    .a(al_1e120105[4]),
    .b(al_1e120105[7]),
    .c(al_1e120105[8]),
    .d(al_2814a16d[4]),
    .e(al_2814a16d[7]),
    .f(al_2814a16d[8]),
    .o(al_e1dab4c9));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_5c5230f5 (
    .a(al_1e120105[0]),
    .b(al_1e120105[5]),
    .c(al_1e120105[10]),
    .d(al_2814a16d[0]),
    .e(al_2814a16d[5]),
    .f(al_2814a16d[10]),
    .o(al_336d8f19));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_c0c4ff24 (
    .a(al_1e120105[6]),
    .b(al_1e120105[9]),
    .c(al_2814a16d[6]),
    .d(al_2814a16d[9]),
    .o(al_9f21cd24));
  AL_MAP_LUT6 #(
    .EQN("~(E*~((D*C*B*A))*~(F)+E*(D*C*B*A)*~(F)+~(E)*(D*C*B*A)*F+E*(D*C*B*A)*F)"),
    .INIT(64'h7fff7fff0000ffff))
    al_5f0fd8ef (
    .a(al_13154bf6),
    .b(al_e1dab4c9),
    .c(al_336d8f19),
    .d(al_9f21cd24),
    .e(al_dacf8588),
    .f(al_e2dc2eea),
    .o(al_b242277f));
  AL_DFF_X al_529a18f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_509509ae),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_dacf8588));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_8206442d (
    .a(al_1a0f7d2b[4]),
    .b(al_1a0f7d2b[5]),
    .c(al_1a0f7d2b[6]),
    .d(al_1a0f7d2b[7]),
    .o(al_162f415f));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*~C*~B*~A)"),
    .INIT(64'h0100000000000000))
    al_10237955 (
    .a(al_74c05d28),
    .b(al_1a0f7d2b[2]),
    .c(al_1a0f7d2b[3]),
    .d(al_b8530805),
    .e(al_fd106601),
    .f(al_ef7f6f7b[1]),
    .o(al_c862ea52));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    al_5f5eafa7 (
    .a(al_c862ea52),
    .b(al_162f415f),
    .c(al_1a0f7d2b[0]),
    .d(al_1a0f7d2b[1]),
    .o(al_ec602117));
  AL_DFF_X al_fc1f1c9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ec602117),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_16c52309));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(C*~(B)*~((E*D))+C*B*~((E*D))+~(C)*B*(E*D)+C*B*(E*D)))"),
    .INIT(32'heefafafa))
    al_2dd9b42b (
    .a(al_6f75ef0e),
    .b(al_1a0f7d2b[0]),
    .c(al_2814a16d[0]),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_13349257[0]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'hfbea))
    al_b513f99c (
    .a(al_6f75ef0e),
    .b(al_ba174b4c),
    .c(al_1a0f7d2b[2]),
    .d(al_2814a16d[10]),
    .o(al_13349257[10]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(C*~(B)*~((E*D))+C*B*~((E*D))+~(C)*B*(E*D)+C*B*(E*D)))"),
    .INIT(32'heefafafa))
    al_49665b12 (
    .a(al_6f75ef0e),
    .b(al_1a0f7d2b[1]),
    .c(al_2814a16d[1]),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_13349257[1]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(C*~(B)*~((E*D))+C*B*~((E*D))+~(C)*B*(E*D)+C*B*(E*D)))"),
    .INIT(32'heefafafa))
    al_e725d714 (
    .a(al_6f75ef0e),
    .b(al_1a0f7d2b[2]),
    .c(al_2814a16d[2]),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_13349257[2]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(C*~(B)*~((E*D))+C*B*~((E*D))+~(C)*B*(E*D)+C*B*(E*D)))"),
    .INIT(32'heefafafa))
    al_55e7cdba (
    .a(al_6f75ef0e),
    .b(al_1a0f7d2b[3]),
    .c(al_2814a16d[3]),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_13349257[3]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(C*~(B)*~((E*D))+C*B*~((E*D))+~(C)*B*(E*D)+C*B*(E*D)))"),
    .INIT(32'heefafafa))
    al_330a3d13 (
    .a(al_6f75ef0e),
    .b(al_1a0f7d2b[4]),
    .c(al_2814a16d[4]),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_13349257[4]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(C*~(B)*~((E*D))+C*B*~((E*D))+~(C)*B*(E*D)+C*B*(E*D)))"),
    .INIT(32'heefafafa))
    al_cc53eb61 (
    .a(al_6f75ef0e),
    .b(al_1a0f7d2b[5]),
    .c(al_2814a16d[5]),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_13349257[5]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(C*~(B)*~((E*D))+C*B*~((E*D))+~(C)*B*(E*D)+C*B*(E*D)))"),
    .INIT(32'heefafafa))
    al_529413a1 (
    .a(al_6f75ef0e),
    .b(al_1a0f7d2b[6]),
    .c(al_2814a16d[6]),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_13349257[6]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(C*~(B)*~((E*D))+C*B*~((E*D))+~(C)*B*(E*D)+C*B*(E*D)))"),
    .INIT(32'heefafafa))
    al_3d682a5a (
    .a(al_6f75ef0e),
    .b(al_1a0f7d2b[7]),
    .c(al_2814a16d[7]),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_13349257[7]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'hfbea))
    al_40a3038 (
    .a(al_6f75ef0e),
    .b(al_ba174b4c),
    .c(al_1a0f7d2b[0]),
    .d(al_2814a16d[8]),
    .o(al_13349257[8]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'hfbea))
    al_e19cf989 (
    .a(al_6f75ef0e),
    .b(al_ba174b4c),
    .c(al_1a0f7d2b[1]),
    .d(al_2814a16d[9]),
    .o(al_13349257[9]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_e3fb7d83 (
    .a(al_162f415f),
    .b(al_1a0f7d2b[0]),
    .c(al_1a0f7d2b[1]),
    .d(al_1a0f7d2b[2]),
    .e(al_1a0f7d2b[3]),
    .o(al_adf11663));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*A)"),
    .INIT(32'h20000000))
    al_b4760851 (
    .a(al_adf11663),
    .b(al_74c05d28),
    .c(al_b8530805),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_d1bf4e26));
  AL_DFF_X al_6b5f8a1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d1bf4e26),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_f9e26d2b));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_bc2edc7a (
    .a(al_adf11663),
    .b(al_ba174b4c),
    .o(al_3fdafe26));
  AL_DFF_X al_4ac5bba (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_3fdafe26),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_b8530805));
  AL_DFF_X al_d5b0e59a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1b7fc148),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_ff7075f1));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    al_c0eeb8c4 (
    .a(al_a409c88e),
    .b(al_4f800f89),
    .c(al_4d5dd241),
    .d(al_ef7f6f7b[0]),
    .o(al_c758ee36));
  AL_MAP_LUT5 #(
    .EQN("((~E*~D*C)*~(B)*~(A)+(~E*~D*C)*B*~(A)+~((~E*~D*C))*B*A+(~E*~D*C)*B*A)"),
    .INIT(32'h888888d8))
    al_f646038f (
    .a(al_c758ee36),
    .b(al_1a0f7d2b[0]),
    .c(al_1b7fc148),
    .d(al_5d14a06f),
    .e(al_bf03de15),
    .o(al_109f9c2b));
  AL_DFF_X al_1f25d7ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_109f9c2b),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1b7fc148));
  AL_DFF_X al_eaba96f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_25af80c5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c3b9f16));
  AL_MAP_LUT6 #(
    .EQN("(~F*~(~A*~(C*~(E*D*B))))"),
    .INIT(64'h00000000bafafafa))
    al_899b6507 (
    .a(al_f9a0f4e),
    .b(rx_clk_en),
    .c(al_8c3b9f16),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .f(al_fea77e50),
    .o(al_25af80c5));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*~C*~B*A)"),
    .INIT(64'h0200000000000000))
    al_1b61a081 (
    .a(rx_clk_en),
    .b(al_1a0f7d2b[6]),
    .c(al_1a0f7d2b[7]),
    .d(al_b8530805),
    .e(al_fd106601),
    .f(al_ef7f6f7b[1]),
    .o(al_96064004));
  AL_MAP_LUT6 #(
    .EQN("(A*~(F*~(~E*~(D*C*B))))"),
    .INIT(64'h00002aaaaaaaaaaa))
    al_934a0824 (
    .a(al_96064004),
    .b(al_1a0f7d2b[1]),
    .c(al_1a0f7d2b[2]),
    .d(al_1a0f7d2b[3]),
    .e(al_1a0f7d2b[4]),
    .f(al_1a0f7d2b[5]),
    .o(al_f9a0f4e));
  AL_DFF_X al_28f542e9 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7ffbbf6e),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ea736991));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_4031331e (
    .a(al_fd106601),
    .b(al_ef7f6f7b[0]),
    .o(al_ba174b4c));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    al_87e0c12e (
    .a(al_162f415f),
    .b(al_1a0f7d2b[1]),
    .c(al_1a0f7d2b[2]),
    .o(al_6f2b16fe));
  AL_MAP_LUT5 #(
    .EQN("~((~E*~B)*~((~D*A))*~(C)+(~E*~B)*(~D*A)*~(C)+~((~E*~B))*(~D*A)*C+(~E*~B)*(~D*A)*C)"),
    .INIT(32'hff5ffc5c))
    al_176d699e (
    .a(al_6f2b16fe),
    .b(al_6f75ef0e),
    .c(al_ba174b4c),
    .d(al_1a0f7d2b[3]),
    .e(al_31cc16da),
    .o(al_29cb9079));
  AL_DFF_X al_ea1efab7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_29cb9079),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_31cc16da));
  AL_DFF_X al_40396ac8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b449eeb9[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_3ccf053a));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_6baca878 (
    .a(al_ba174b4c),
    .b(al_1a0f7d2b[4]),
    .c(al_1a0f7d2b[5]),
    .d(al_1a0f7d2b[6]),
    .e(al_1a0f7d2b[7]),
    .o(al_4c3c2401));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*C*B*A)"),
    .INIT(64'h0000000000000080))
    al_96014cb0 (
    .a(al_4c3c2401),
    .b(al_e646046),
    .c(al_1a0f7d2b[0]),
    .d(al_1a0f7d2b[1]),
    .e(al_1a0f7d2b[2]),
    .f(al_1a0f7d2b[3]),
    .o(al_f97fd11e));
  AL_MAP_LUT6 #(
    .EQN("((~D*C)*~((B*A))*~((F*E))+(~D*C)*(B*A)*~((F*E))+~((~D*C))*(B*A)*(F*E)+(~D*C)*(B*A)*(F*E))"),
    .INIT(64'h888800f000f000f0))
    al_97b7d3a3 (
    .a(al_adf11663),
    .b(al_b449eeb9[0]),
    .c(al_b449eeb9[1]),
    .d(al_5d14a06f),
    .e(al_fd106601),
    .f(al_ef7f6f7b[1]),
    .o(al_46118f46));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_bc03f167 (
    .a(1'b0),
    .o({al_95894036,open_n6}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_29d9ad55 (
    .a(al_b9d3b2c1[0]),
    .b(1'b1),
    .c(al_95894036),
    .o({al_6fed1e72,al_66bdfa10[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_507e1816 (
    .a(al_b9d3b2c1[1]),
    .b(1'b0),
    .c(al_6fed1e72),
    .o({al_8f867af4,al_66bdfa10[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d1e6557b (
    .a(al_b9d3b2c1[2]),
    .b(1'b0),
    .c(al_8f867af4),
    .o({al_f03499fc,al_66bdfa10[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5031517c (
    .a(al_b9d3b2c1[3]),
    .b(1'b0),
    .c(al_f03499fc),
    .o({al_db3e7a3b,al_66bdfa10[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1953411a (
    .a(al_b9d3b2c1[4]),
    .b(1'b0),
    .c(al_db3e7a3b),
    .o({al_f1799bbf,al_66bdfa10[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b5d16cce (
    .a(al_b9d3b2c1[5]),
    .b(1'b0),
    .c(al_f1799bbf),
    .o({al_c5cae25a,al_66bdfa10[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a4d4e3f8 (
    .a(al_b9d3b2c1[6]),
    .b(1'b0),
    .c(al_c5cae25a),
    .o({al_6f517dcb,al_66bdfa10[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_93d8792e (
    .a(al_b9d3b2c1[7]),
    .b(1'b0),
    .c(al_6f517dcb),
    .o({al_5d55f7bd,al_66bdfa10[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_60faeef3 (
    .a(al_b9d3b2c1[8]),
    .b(1'b0),
    .c(al_5d55f7bd),
    .o({al_93f12ca5,al_66bdfa10[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3d2e3998 (
    .a(al_b9d3b2c1[9]),
    .b(1'b0),
    .c(al_93f12ca5),
    .o({al_822d50d7,al_66bdfa10[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3becfa36 (
    .a(al_b9d3b2c1[10]),
    .b(1'b0),
    .c(al_822d50d7),
    .o({al_be626253,al_66bdfa10[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3f2bd598 (
    .a(al_b9d3b2c1[11]),
    .b(1'b0),
    .c(al_be626253),
    .o({al_55aaf816,al_66bdfa10[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cdc2510b (
    .a(al_b9d3b2c1[12]),
    .b(1'b0),
    .c(al_55aaf816),
    .o({al_a5f70472,al_66bdfa10[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4773d331 (
    .a(al_b9d3b2c1[13]),
    .b(1'b0),
    .c(al_a5f70472),
    .o({al_5c2a2da8,al_66bdfa10[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3ab12c1f (
    .a(al_b9d3b2c1[14]),
    .b(1'b0),
    .c(al_5c2a2da8),
    .o({open_n7,al_66bdfa10[14]}));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_9aadf015 (
    .a(rx_clk_en),
    .b(al_ea736991),
    .c(al_b9d3b2c1[14]),
    .o(al_65f65cdd));
  AL_DFF_X al_dd4b9270 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[8]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[8]));
  AL_DFF_X al_cc286e64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[9]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[9]));
  AL_DFF_X al_ab0120e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[10]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[10]));
  AL_DFF_X al_b1a00dbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[0]));
  AL_DFF_X al_728ed1f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[1]));
  AL_DFF_X al_9520b60e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[2]));
  AL_DFF_X al_74a75b7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[3]));
  AL_DFF_X al_9b82cfda (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[4]));
  AL_DFF_X al_201de3fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[5]));
  AL_DFF_X al_fc2e09f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[6]));
  AL_DFF_X al_42668359 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ea827a0c[7]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1e120105[7]));
  AL_DFF_X al_57caed84 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[8]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[8]));
  AL_DFF_X al_d52d3752 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[9]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[9]));
  AL_DFF_X al_23febcf2 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[10]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[10]));
  AL_DFF_X al_b700ad3c (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[11]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[11]));
  AL_DFF_X al_2546face (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[12]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[12]));
  AL_DFF_X al_5b82fa1b (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[13]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[13]));
  AL_DFF_X al_381ea887 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[14]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[14]));
  AL_DFF_X al_3b888006 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[0]));
  AL_DFF_X al_80984e (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[1]));
  AL_DFF_X al_d45489ad (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[2]));
  AL_DFF_X al_3fa0bc7e (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[3]));
  AL_DFF_X al_53a7f8b9 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[4]));
  AL_DFF_X al_89f39c4a (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[5]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[5]));
  AL_DFF_X al_7bc0c667 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[6]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[6]));
  AL_DFF_X al_4150cc3f (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e843f7[7]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9d3b2c1[7]));
  AL_DFF_X al_984b19d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[8]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[8]));
  AL_DFF_X al_7c5f6570 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[9]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[9]));
  AL_DFF_X al_a259ad7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[10]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[10]));
  AL_DFF_X al_f917a9c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[0]));
  AL_DFF_X al_c452fb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[1]));
  AL_DFF_X al_37be32c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[2]));
  AL_DFF_X al_de90691 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[3]));
  AL_DFF_X al_443655a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[4]));
  AL_DFF_X al_c7dc10a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[5]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[5]));
  AL_DFF_X al_3bb18f78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[6]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[6]));
  AL_DFF_X al_210820b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_13349257[7]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_2814a16d[7]));
  AL_DFF_X al_7fe39dd9 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[8]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[8]));
  AL_DFF_X al_3fe03c5c (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[9]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[9]));
  AL_DFF_X al_2ad8f411 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[10]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[10]));
  AL_DFF_X al_626a58a5 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[11]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[11]));
  AL_DFF_X al_a66bfd41 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[12]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[12]));
  AL_DFF_X al_89ec3eca (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[13]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[13]));
  AL_DFF_X al_31b236d1 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[0]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[0]));
  AL_DFF_X al_1dafad22 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[1]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[1]));
  AL_DFF_X al_2f63bb62 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[2]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[2]));
  AL_DFF_X al_3e3a2a19 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[3]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[3]));
  AL_DFF_X al_99ebaa8 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[4]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[4]));
  AL_DFF_X al_3df4efb4 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[5]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[5]));
  AL_DFF_X al_b8f88af6 (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[6]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[6]));
  AL_DFF_X al_b117def (
    .ar(al_fea77e50),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9d3b2c1[7]),
    .en(al_65f65cdd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26b248e8[7]));
  AL_DFF_X al_d8dbe81f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f97fd11e),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_b449eeb9[0]));
  AL_DFF_X al_b5e34de7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_46118f46),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_b449eeb9[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_cbcd5e30 (
    .a(al_cc7e79c9),
    .b(al_d6bd6336),
    .o(al_82dda9be));
  AL_DFF_X al_b90bbaea (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_82dda9be),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_c99d4c23));
  AL_DFF_X al_b28afc55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b8f86eed),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9cabf6c6));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*~(C)*~((B*A))+D*C*~((B*A))+~(D)*C*(B*A)+D*C*(B*A)))"),
    .INIT(32'hfffff780))
    al_d9581e80 (
    .a(al_153d6f9e),
    .b(rx_clk_en),
    .c(al_677d00f0[2]),
    .d(al_9cabf6c6),
    .e(al_fea77e50),
    .o(al_b8f86eed));
  AL_DFF_X al_50b78e3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_597cc1f6),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_b19043fc));
  AL_DFF_X al_4d7e4915 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b0b9c021),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_225d06ad));
  AL_MAP_LUT5 #(
    .EQN("(~E*(D*~(C)*~((B*A))+D*C*~((B*A))+~(D)*C*(B*A)+D*C*(B*A)))"),
    .INIT(32'h0000f780))
    al_5513850f (
    .a(al_6f75ef0e),
    .b(rx_clk_en),
    .c(al_677d00f0[5]),
    .d(al_225d06ad),
    .e(al_fea77e50),
    .o(al_b0b9c021));
  AL_DFF_X al_856afeda (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8cebb59e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_74c05d28));
  AL_MAP_LUT5 #(
    .EQN("(~E*(D*~(C)*~((B*A))+D*C*~((B*A))+~(D)*C*(B*A)+D*C*(B*A)))"),
    .INIT(32'h0000f780))
    al_720817c3 (
    .a(al_6f75ef0e),
    .b(rx_clk_en),
    .c(al_677d00f0[6]),
    .d(al_74c05d28),
    .e(al_fea77e50),
    .o(al_8cebb59e));
  AL_DFF_X al_316e57af (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4ab032f9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6d3d88));
  AL_MAP_LUT5 #(
    .EQN("(~E*(D*~(C)*~((B*A))+D*C*~((B*A))+~(D)*C*(B*A)+D*C*(B*A)))"),
    .INIT(32'h0000f780))
    al_3d31c830 (
    .a(al_6f75ef0e),
    .b(rx_clk_en),
    .c(al_677d00f0[7]),
    .d(al_6c6d3d88),
    .e(al_fea77e50),
    .o(al_4ab032f9));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_1f1c5811 (
    .a(al_e729b3e2),
    .b(al_6133949d[3]),
    .c(al_bd413a73[3]),
    .d(al_e799d30a[3]),
    .o(al_597cc1f6));
  AL_DFF_X al_e60b793 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_16302c3d),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_d83e61fb));
  AL_DFF_X al_6aee0ed7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d83e61fb),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_932a07c7));
  AL_DFF_X al_d894dbd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_469f2a04[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_62730356));
  AL_DFF_X al_90c4e8f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_62730356),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7ffbbf6e));
  AL_DFF_X al_6b77e12f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_60057698),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7a7628f9));
  AL_DFF_X al_2e5b6757 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ff43a01c[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_ebdfe328));
  AL_DFF_X al_c03a4dd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ebdfe328),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7c1aee64));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(~C*A))"),
    .INIT(8'hce))
    al_544f6a1e (
    .a(al_a409c88e),
    .b(al_4d5dd241),
    .c(al_2c3ff84c),
    .o(al_4360005c));
  AL_DFF_X al_765c4df4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4360005c),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_a409c88e));
  AL_MAP_LUT5 #(
    .EQN("(~C*A*~(~B*~(E*D)))"),
    .INIT(32'h0a080808))
    al_60bd08df (
    .a(al_62730356),
    .b(al_e2dc2eea),
    .c(al_4d5dd241),
    .d(al_fd106601),
    .e(al_ef7f6f7b[1]),
    .o(al_f0362cc));
  AL_DFF_X al_9180c5e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0362cc),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_e2dc2eea));
  AL_MAP_LUT6 #(
    .EQN("(~F*A*~(~D*~(C*~(~E*B))))"),
    .INIT(64'h00000000aaa0aa20))
    al_3d313cdb (
    .a(al_62730356),
    .b(al_7ffbbf6e),
    .c(al_cb67e17c),
    .d(al_4f800f89),
    .e(al_db678397),
    .f(al_ef7f6f7b[5]),
    .o(al_d5a6be8d));
  AL_DFF_X al_33c508c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d5a6be8d),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_4f800f89));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_825d2d39 (
    .a(al_d83e61fb),
    .b(al_932a07c7),
    .o(al_ce94a07b));
  AL_DFF_X al_17fcb203 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ce94a07b),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_4d5dd241));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_93b97c0 (
    .a(al_e729b3e2),
    .b(al_6133949d[3]),
    .c(al_bd413a73[3]),
    .d(al_e799d30a[3]),
    .o(al_9809ce8b));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~(C*~B*~A))"),
    .INIT(32'h00ef0000))
    al_2998ee35 (
    .a(al_9809ce8b),
    .b(al_469f2a04[2]),
    .c(al_ff43a01c[3]),
    .d(al_6598ce3a),
    .e(al_8fc9814c),
    .o(al_9e79b57b));
  AL_DFF_X al_f24645d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9e79b57b),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_6598ce3a));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_83b8c397 (
    .a(al_62730356),
    .b(al_469f2a04[2]),
    .o(al_b1f059e9));
  AL_DFF_X al_9ce36048 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b1f059e9),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_2c3ff84c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*~A)"),
    .INIT(64'h0000000000000004))
    al_955842e8 (
    .a(al_469f2a04[2]),
    .b(al_ff43a01c[3]),
    .c(al_ddf438c2[3]),
    .d(al_33bfe5eb[3]),
    .e(al_dd83fb37[3]),
    .f(al_7bd9ce9a[3]),
    .o(al_9b66e5cd));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9805d0c3 (
    .a(al_9b66e5cd),
    .b(al_4c32576a[3]),
    .o(al_e729b3e2));
  AL_MAP_LUT6 #(
    .EQN("(~C*B*~(A*(~(D)*~(E)*~(F)+D*E*F)))"),
    .INIT(64'h040c0c0c0c0c0c04))
    al_cbddb182 (
    .a(al_e729b3e2),
    .b(al_ebdfe328),
    .c(al_f02638e3),
    .d(al_6133949d[3]),
    .e(al_bd413a73[3]),
    .f(al_e799d30a[3]),
    .o(al_9f6030e));
  AL_MAP_LUT6 #(
    .EQN("(~F*~D*~(~E*~(C*~B*~A)))"),
    .INIT(64'h0000000000ff0010))
    al_3db725c4 (
    .a(al_7ffbbf6e),
    .b(al_ebdfe328),
    .c(al_7c1aee64),
    .d(al_f02638e3),
    .e(al_6598ce3a),
    .f(al_5d14a06f),
    .o(al_b9b188f3));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D*~C*~A))"),
    .INIT(16'hcdcc))
    al_ca9bfbae (
    .a(al_9f6030e),
    .b(al_b9b188f3),
    .c(al_62730356),
    .d(al_7ffbbf6e),
    .o(al_debb55eb));
  AL_DFF_X al_85523685 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_debb55eb),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5d14a06f));
  AL_MAP_LUT6 #(
    .EQN("(D*~C*~B*~A*~(~F*~E))"),
    .INIT(64'h0100010001000000))
    al_8ad50a2c (
    .a(al_6e672ebc),
    .b(al_b19043fc),
    .c(al_62730356),
    .d(al_ebdfe328),
    .e(al_a409c88e),
    .f(al_8fc9814c),
    .o(al_50559550));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_675e6c91 (
    .a(al_50559550),
    .b(al_f02638e3),
    .o(al_b99dff45));
  AL_DFF_X al_fd6ad9ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b99dff45),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_8fc9814c));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_ebac1e95 (
    .a(al_5d14a06f),
    .b(al_ef7f6f7b[1]),
    .o(al_6aa6d3c8[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_7f6a83c4 (
    .a(al_5d14a06f),
    .b(al_ef7f6f7b[2]),
    .o(al_6aa6d3c8[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_42473f89 (
    .a(al_5d14a06f),
    .b(al_ef7f6f7b[3]),
    .o(al_6aa6d3c8[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_8eaf14be (
    .a(al_5d14a06f),
    .b(al_ef7f6f7b[4]),
    .o(al_6aa6d3c8[3]));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~C*~(~E*~D*~B*~A))"),
    .INIT(64'hfffffffff0f0f0f1))
    al_cf8c795d (
    .a(al_a409c88e),
    .b(al_4f800f89),
    .c(al_5d14a06f),
    .d(al_fd106601),
    .e(al_5b221454),
    .f(al_ef7f6f7b[5]),
    .o(al_4ceb8d18[0]));
  AL_MAP_LUT6 #(
    .EQN("(F*~C*~(~E*~D*~B*~A))"),
    .INIT(64'h0f0f0f0e00000000))
    al_1be4d24c (
    .a(al_a409c88e),
    .b(al_4f800f89),
    .c(al_5d14a06f),
    .d(al_fd106601),
    .e(al_5b221454),
    .f(al_ef7f6f7b[0]),
    .o(al_4ceb8d18[1]));
  AL_MAP_LUT5 #(
    .EQN("(~D*A*~(~B*~(E*C)))"),
    .INIT(32'h00a80088))
    al_69aff296 (
    .a(al_62730356),
    .b(al_fd106601),
    .c(al_5b221454),
    .d(al_ef7f6f7b[1]),
    .e(al_ef7f6f7b[5]),
    .o(al_ca4883db));
  AL_DFF_X al_138df406 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ca4883db),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_fd106601));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~(E*~D)*~(~C*A)))"),
    .INIT(32'h08cc0808))
    al_ed1487e2 (
    .a(al_4c9b2533),
    .b(al_62730356),
    .c(al_7ffbbf6e),
    .d(al_cb67e17c),
    .e(al_db678397),
    .o(al_cb7ab50c));
  AL_DFF_X al_42c1556a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cb7ab50c),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_db678397));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h88a0))
    al_e4146969 (
    .a(al_62730356),
    .b(al_4f800f89),
    .c(al_5b221454),
    .d(al_ef7f6f7b[5]),
    .o(al_53cf6c8d));
  AL_DFF_X al_11e38a47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53cf6c8d),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5b221454));
  AL_DFF_X al_8a35e174 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4ceb8d18[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_fea77e50),
    .q(al_ef7f6f7b[0]));
  AL_DFF_X al_77998ea7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4ceb8d18[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_ef7f6f7b[1]));
  AL_DFF_X al_2a2fc392 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6aa6d3c8[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_ef7f6f7b[2]));
  AL_DFF_X al_4dd19fe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6aa6d3c8[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_ef7f6f7b[3]));
  AL_DFF_X al_a0ba4d4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6aa6d3c8[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_ef7f6f7b[4]));
  AL_DFF_X al_1c39c0c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6aa6d3c8[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_ef7f6f7b[5]));
  AL_DFF_X al_f38b8fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_48908c7b),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vld));
  AL_MAP_LUT6 #(
    .EQN("(F*E*~D*C*~B*A)"),
    .INIT(64'h0020000000000000))
    al_c573dc13 (
    .a(al_1d03242c[2]),
    .b(al_1d03242c[3]),
    .c(al_1d03242c[4]),
    .d(al_1d03242c[5]),
    .e(al_1d03242c[6]),
    .f(al_1d03242c[7]),
    .o(al_4e1502ae));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    al_27f35f01 (
    .a(al_4e1502ae),
    .b(al_62730356),
    .c(al_ebdfe328),
    .d(al_1d03242c[0]),
    .e(al_1d03242c[1]),
    .o(al_5274ea30));
  AL_DFF_X al_9a97493b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5274ea30),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_cb67e17c));
  AL_DFF_X al_d0b247b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_72bd37a4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f02638e3));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~D*~(C)*~((B*A))+~D*C*~((B*A))+~(~D)*C*(B*A)+~D*C*(B*A)))"),
    .INIT(32'h00007f08))
    al_2eccffea (
    .a(al_6f75ef0e),
    .b(rx_clk_en),
    .c(al_44560df6[1]),
    .d(al_f02638e3),
    .e(al_fea77e50),
    .o(al_72bd37a4));
  AL_DFF_X al_82b19848 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_60b3be17),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_48908c7b));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d963cc5a (
    .a(al_18642257),
    .b(al_e5a67968),
    .o(al_54280ae3[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_61a9c62a (
    .a(al_18642257),
    .b(al_e5a67968),
    .o(al_54280ae3[1]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_619a863b (
    .a(al_a6104abc),
    .b(al_a3910e3c),
    .o(al_4c1d19df));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*~(~B*~(E*A)))"),
    .INIT(32'h000e000c))
    al_30bd88ff (
    .a(al_4c1d19df),
    .b(al_cc7e79c9),
    .c(al_e1057698),
    .d(al_d6bd6336),
    .e(al_7ac96e46),
    .o(al_91fb7c78));
  AL_DFF_X al_9396d50a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_91fb7c78),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_cc7e79c9));
  AL_DFF_X al_7e18da5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b2e646bb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e646046));
  AL_MAP_LUT5 #(
    .EQN("(~E*(D*~(C)*~((B*A))+D*C*~((B*A))+~(D)*C*(B*A)+D*C*(B*A)))"),
    .INIT(32'h0000f780))
    al_4e36ea7c (
    .a(al_6f75ef0e),
    .b(rx_clk_en),
    .c(al_677d00f0[3]),
    .d(al_e646046),
    .e(al_fea77e50),
    .o(al_b2e646bb));
  AL_DFF_X al_57112a5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5e036bbd[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_aeb75558[0]));
  AL_DFF_X al_46edc48b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5e036bbd[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_aeb75558[1]));
  AL_DFF_X al_dcc940e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5e036bbd[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_aeb75558[2]));
  AL_DFF_X al_1a6606af (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5e036bbd[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_aeb75558[3]));
  AL_DFF_X al_c4d7fb66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5e036bbd[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_aeb75558[4]));
  AL_DFF_X al_fb7973fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5e036bbd[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_aeb75558[5]));
  AL_DFF_X al_e0767e34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5e036bbd[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_aeb75558[6]));
  AL_DFF_X al_f499aa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5e036bbd[7]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_aeb75558[7]));
  AL_DFF_X al_a8c067ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53486c5d[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_583c216b[0]));
  AL_DFF_X al_3e53d8c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53486c5d[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_583c216b[1]));
  AL_DFF_X al_7c74f893 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53486c5d[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_583c216b[2]));
  AL_DFF_X al_bd70c39c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53486c5d[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_583c216b[3]));
  AL_DFF_X al_97603391 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53486c5d[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_583c216b[4]));
  AL_DFF_X al_d6dff8be (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53486c5d[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_583c216b[5]));
  AL_DFF_X al_95be80ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53486c5d[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_583c216b[6]));
  AL_DFF_X al_1f292a10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53486c5d[7]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_583c216b[7]));
  AL_DFF_X al_3e9a2558 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ddf438c2[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1d03242c[0]));
  AL_DFF_X al_ae52895d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6133949d[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1d03242c[1]));
  AL_DFF_X al_1a478332 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_bd413a73[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1d03242c[2]));
  AL_DFF_X al_67a5c15b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e799d30a[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1d03242c[3]));
  AL_DFF_X al_5b89d103 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_33bfe5eb[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1d03242c[4]));
  AL_DFF_X al_a50c2432 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_dd83fb37[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1d03242c[5]));
  AL_DFF_X al_7dbb340e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7bd9ce9a[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1d03242c[6]));
  AL_DFF_X al_6d830c6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4c32576a[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1d03242c[7]));
  AL_DFF_X al_f5953ee0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1d03242c[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1a0f7d2b[0]));
  AL_DFF_X al_953fbfa0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1d03242c[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1a0f7d2b[1]));
  AL_DFF_X al_e43b3f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1d03242c[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1a0f7d2b[2]));
  AL_DFF_X al_9a586125 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1d03242c[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1a0f7d2b[3]));
  AL_DFF_X al_ec6a2fa9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1d03242c[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1a0f7d2b[4]));
  AL_DFF_X al_41ff88fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1d03242c[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1a0f7d2b[5]));
  AL_DFF_X al_1720861d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1d03242c[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1a0f7d2b[6]));
  AL_DFF_X al_44f43963 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1d03242c[7]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_1a0f7d2b[7]));
  AL_DFF_X al_10c0f018 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1a0f7d2b[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5e036bbd[0]));
  AL_DFF_X al_8749ee34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1a0f7d2b[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5e036bbd[1]));
  AL_DFF_X al_5f916498 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1a0f7d2b[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5e036bbd[2]));
  AL_DFF_X al_84245345 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1a0f7d2b[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5e036bbd[3]));
  AL_DFF_X al_1ef04064 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1a0f7d2b[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5e036bbd[4]));
  AL_DFF_X al_f91ed01c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1a0f7d2b[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5e036bbd[5]));
  AL_DFF_X al_e2985245 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1a0f7d2b[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5e036bbd[6]));
  AL_DFF_X al_bfe5be51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1a0f7d2b[7]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5e036bbd[7]));
  AL_DFF_X al_169e5e33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[8]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[8]));
  AL_DFF_X al_1b7f0140 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[9]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[9]));
  AL_DFF_X al_2b4fa843 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[10]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[10]));
  AL_DFF_X al_c35f6b76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[11]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[11]));
  AL_DFF_X al_271b5296 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[12]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[12]));
  AL_DFF_X al_ea7da777 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[13]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[13]));
  AL_DFF_X al_ce389adf (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[14]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[14]));
  AL_DFF_X al_498005f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[15]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[15]));
  AL_DFF_X al_9af14e91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[16]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[16]));
  AL_DFF_X al_90ba25c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[17]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[17]));
  AL_DFF_X al_11be304b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[0]));
  AL_DFF_X al_aa59c4a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[18]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[18]));
  AL_DFF_X al_c4eb13f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[19]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[21]));
  AL_DFF_X al_59ac8051 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[20]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[19]));
  AL_DFF_X al_e661489b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[21]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[22]));
  AL_DFF_X al_ffcd1d0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[23]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[20]));
  AL_DFF_X al_285625d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[24]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[25]));
  AL_DFF_X al_159561bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[1]));
  AL_DFF_X al_71197b2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[26]));
  AL_DFF_X al_1febb41e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[2]));
  AL_DFF_X al_851b0725 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[3]));
  AL_DFF_X al_eba1611 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[5]));
  AL_DFF_X al_6820bada (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[6]));
  AL_DFF_X al_c4a953e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_36654522[7]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[7]));
  AL_DFF_X al_1e8eb3bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[8]));
  AL_DFF_X al_1327679d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[4]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[9]));
  AL_DFF_X al_dcc81112 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[10]));
  AL_DFF_X al_7ed91db5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[6]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[11]));
  AL_DFF_X al_b9feef6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[7]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[12]));
  AL_DFF_X al_d93d7fc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[8]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[13]));
  AL_DFF_X al_1f7a6b72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[9]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[14]));
  AL_DFF_X al_6916559a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[10]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[15]));
  AL_DFF_X al_639a4d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[11]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[16]));
  AL_DFF_X al_b496d0a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[12]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[17]));
  AL_DFF_X al_26eb3239 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d6bd6336),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[0]));
  AL_DFF_X al_fcf9c4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[13]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[18]));
  AL_DFF_X al_c02a1c40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ce99d34),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[19]));
  AL_DFF_X al_7f15cecb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f5080327),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[20]));
  AL_DFF_X al_4885de2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_3ccf053a),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[21]));
  AL_DFF_X al_224b57d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b95885c7),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[23]));
  AL_DFF_X al_ac906732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_54280ae3[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[24]));
  AL_DFF_X al_85a88830 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1057698),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[1]));
  AL_DFF_X al_ba74bbb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_54280ae3[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[2]));
  AL_DFF_X al_ee1183a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_81b839ee[5]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[3]));
  AL_DFF_X al_52303269 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ff7075f1),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[4]));
  AL_DFF_X al_e13d4617 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[5]));
  AL_DFF_X al_9e8b7a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[6]));
  AL_DFF_X al_c3957944 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_26b248e8[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_36654522[7]));
  AL_DFF_0 al_bd59e6ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_583c216b[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ddf438c2[0]));
  AL_DFF_0 al_48e2644e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ddf438c2[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ddf438c2[1]));
  AL_DFF_0 al_474d1336 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ddf438c2[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ddf438c2[2]));
  AL_DFF_0 al_b3489d3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ddf438c2[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ddf438c2[3]));
  AL_DFF_0 al_4a5d2335 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_583c216b[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6133949d[0]));
  AL_DFF_0 al_b86ce009 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6133949d[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6133949d[1]));
  AL_DFF_0 al_4427a7be (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6133949d[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6133949d[2]));
  AL_DFF_0 al_e7d8bd2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6133949d[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6133949d[3]));
  AL_DFF_0 al_c3b954ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_583c216b[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd413a73[0]));
  AL_DFF_0 al_d842ce34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_bd413a73[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd413a73[1]));
  AL_DFF_0 al_17ed2f1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_bd413a73[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd413a73[2]));
  AL_DFF_0 al_69233b59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_bd413a73[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd413a73[3]));
  AL_DFF_0 al_7d86f9f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_583c216b[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e799d30a[0]));
  AL_DFF_0 al_6609820e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e799d30a[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e799d30a[1]));
  AL_DFF_0 al_be6f3d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e799d30a[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e799d30a[2]));
  AL_DFF_0 al_6606d074 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e799d30a[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e799d30a[3]));
  AL_DFF_0 al_c020f3b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_583c216b[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33bfe5eb[0]));
  AL_DFF_0 al_b3cdbb06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_33bfe5eb[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33bfe5eb[1]));
  AL_DFF_0 al_71e55241 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_33bfe5eb[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33bfe5eb[2]));
  AL_DFF_0 al_fbc36806 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_33bfe5eb[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33bfe5eb[3]));
  AL_DFF_0 al_dfa5981d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_583c216b[5]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd83fb37[0]));
  AL_DFF_0 al_8afd8438 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_dd83fb37[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd83fb37[1]));
  AL_DFF_0 al_9f7476ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_dd83fb37[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd83fb37[2]));
  AL_DFF_0 al_3f135b7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_dd83fb37[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd83fb37[3]));
  AL_DFF_0 al_a474c78d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_583c216b[6]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7bd9ce9a[0]));
  AL_DFF_0 al_5c18029 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7bd9ce9a[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7bd9ce9a[1]));
  AL_DFF_0 al_6fb5c22f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7bd9ce9a[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7bd9ce9a[2]));
  AL_DFF_0 al_abf9d478 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7bd9ce9a[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7bd9ce9a[3]));
  AL_DFF_0 al_f763e17d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_583c216b[7]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c32576a[0]));
  AL_DFF_0 al_244ef03d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4c32576a[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c32576a[1]));
  AL_DFF_0 al_f8c67a23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4c32576a[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c32576a[2]));
  AL_DFF_0 al_1ff91315 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4c32576a[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c32576a[3]));
  AL_DFF_X al_37aec6c3 (
    .ar(1'b0),
    .as(al_156e79c6),
    .clk(rx_mac_clk),
    .d(1'b0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d123240));
  AL_DFF_X al_24cd6944 (
    .ar(1'b0),
    .as(al_156e79c6),
    .clk(rx_mac_clk),
    .d(al_7d123240),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_58a58247));
  AL_DFF_X al_c3a92415 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_58a58247),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_379fd30a));
  AL_DFF_X al_1ec58119 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_72818778),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fea77e50));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_272b11c7 (
    .a(al_58a58247),
    .b(al_379fd30a),
    .o(al_72818778));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_1d035f72 (
    .a(reset),
    .b(al_677d00f0[0]),
    .o(al_156e79c6));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9dab6803 (
    .a(al_44560df6[0]),
    .b(al_44560df6[1]),
    .o(al_e48259f9));
  AL_DFF_0 al_f00bcf57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_e48259f9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(speed_100));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_a6064aa9 (
    .a(al_44560df6[1]),
    .o(al_7b681f71));
  AL_DFF_0 al_33366491 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7b681f71),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b821ca29));
  AL_DFF_X al_e4758f02 (
    .ar(1'b0),
    .as(al_aff8bba6),
    .clk(tx_mac_clk),
    .d(1'b0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ceee241e));
  AL_DFF_X al_73d5fb7b (
    .ar(1'b0),
    .as(al_aff8bba6),
    .clk(tx_mac_clk),
    .d(al_ceee241e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a71f4bd6));
  AL_DFF_X al_75d028a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a71f4bd6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a296c440));
  AL_DFF_X al_4e8a3693 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9fbc578a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2dbca608));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_1010a256 (
    .a(al_a71f4bd6),
    .b(al_a296c440),
    .o(al_9fbc578a));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_b2981168 (
    .a(reset),
    .b(al_32c99495[0]),
    .o(al_aff8bba6));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_374d481e (
    .a(al_c9168fb8[3]),
    .o(al_21330e1d[1]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_66fe83f6 (
    .a(al_c9168fb8[4]),
    .o(al_21330e1d[2]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_197e038b (
    .a(al_c9168fb8[5]),
    .o(al_21330e1d[3]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_5e2d640d (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[0]),
    .d(al_90205973[1]),
    .o(al_69384d3c[0]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_d8b197a3 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[10]),
    .d(al_90205973[11]),
    .o(al_69384d3c[10]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_86a4a523 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[11]),
    .d(al_90205973[12]),
    .o(al_69384d3c[11]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_6fbe5d20 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[12]),
    .d(al_90205973[13]),
    .o(al_69384d3c[12]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_bee6119f (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[13]),
    .d(al_90205973[14]),
    .o(al_69384d3c[13]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_a701689 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[1]),
    .d(al_90205973[2]),
    .o(al_69384d3c[1]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_d4445927 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[2]),
    .d(al_90205973[3]),
    .o(al_69384d3c[2]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_75971ee1 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[3]),
    .d(al_90205973[4]),
    .o(al_69384d3c[3]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_83e0d9e (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[4]),
    .d(al_90205973[5]),
    .o(al_69384d3c[4]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_81b9c8c2 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[5]),
    .d(al_90205973[6]),
    .o(al_69384d3c[5]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_fa38d4eb (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[6]),
    .d(al_90205973[7]),
    .o(al_69384d3c[6]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_dd5694cb (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[7]),
    .d(al_90205973[8]),
    .o(al_69384d3c[7]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_be175944 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[8]),
    .d(al_90205973[9]),
    .o(al_69384d3c[8]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_dd216a82 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_90205973[9]),
    .d(al_90205973[10]),
    .o(al_69384d3c[9]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_262df5cc (
    .a(al_90205973[13]),
    .b(al_90205973[14]),
    .o(al_95293982));
  AL_DFF_X al_5595ed8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[8]));
  AL_DFF_X al_31ad334 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[9]));
  AL_DFF_X al_253ae86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[10]));
  AL_DFF_X al_bf1c8ddb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[11]));
  AL_DFF_X al_50d0d252 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[12]));
  AL_DFF_X al_76bd3267 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[13]));
  AL_DFF_X al_4e4debf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[14]));
  AL_DFF_X al_c422ade4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_95293982),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_90205973[0]));
  AL_DFF_X al_2e5cdc19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[1]));
  AL_DFF_X al_46a1e6dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[2]));
  AL_DFF_X al_6982f06c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[3]));
  AL_DFF_X al_562eb7df (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[4]));
  AL_DFF_X al_92ccde50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[5]));
  AL_DFF_X al_2512c3dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[6]));
  AL_DFF_X al_4233808b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_69384d3c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90205973[7]));
  AL_DFF_X al_2c16525d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa981a62[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aa981a62[8]));
  AL_DFF_X al_e6024c7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa981a62[8]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aa981a62[9]));
  AL_DFF_X al_7612488c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_90205973[14]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aa981a62[0]));
  AL_DFF_X al_8e06a4cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa981a62[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aa981a62[1]));
  AL_DFF_X al_2539c511 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa981a62[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aa981a62[2]));
  AL_DFF_X al_4a5d533f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa981a62[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aa981a62[3]));
  AL_DFF_X al_ad59480a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa981a62[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aa981a62[4]));
  AL_DFF_X al_6738f0ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa981a62[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aa981a62[5]));
  AL_DFF_X al_cb814e1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa981a62[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aa981a62[6]));
  AL_DFF_X al_37aa5627 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa981a62[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aa981a62[7]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(~D*~C*B))"),
    .INIT(16'h555d))
    al_23d9495d (
    .a(al_a21ad81c[0]),
    .b(al_fff0fd72[0]),
    .c(al_fff0fd72[1]),
    .d(al_fff0fd72[2]),
    .o(al_acfeaf96[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~D*C)*~(B@A))"),
    .INIT(32'h99999909))
    al_eca4cae2 (
    .a(al_a21ad81c[0]),
    .b(al_a21ad81c[1]),
    .c(al_fff0fd72[0]),
    .d(al_fff0fd72[1]),
    .e(al_fff0fd72[2]),
    .o(al_acfeaf96[1]));
  AL_MAP_LUT6 #(
    .EQN("~(~(~F*~E*D)*~(C@(~B*~A)))"),
    .INIT(64'he1e1e1e1e1e1ffe1))
    al_2c068e49 (
    .a(al_a21ad81c[0]),
    .b(al_a21ad81c[1]),
    .c(al_a21ad81c[2]),
    .d(al_fff0fd72[0]),
    .e(al_fff0fd72[1]),
    .f(al_fff0fd72[2]),
    .o(al_acfeaf96[2]));
  AL_MAP_LUT4 #(
    .EQN("(D@(~C*~B*~A))"),
    .INIT(16'hfe01))
    al_43a52e80 (
    .a(al_a21ad81c[0]),
    .b(al_a21ad81c[1]),
    .c(al_a21ad81c[2]),
    .d(al_a21ad81c[3]),
    .o(al_64a47488[3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*B))"),
    .INIT(16'haaa2))
    al_8178bfaa (
    .a(al_64a47488[3]),
    .b(al_fff0fd72[0]),
    .c(al_fff0fd72[1]),
    .d(al_fff0fd72[2]),
    .o(al_acfeaf96[3]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(C)*~((~D*~B*~A))+E*C*~((~D*~B*~A))+~(E)*C*(~D*~B*~A)+E*C*(~D*~B*~A))"),
    .INIT(32'hfffe0010))
    al_cbbc0b56 (
    .a(al_a21ad81c[0]),
    .b(al_a21ad81c[1]),
    .c(al_a21ad81c[2]),
    .d(al_a21ad81c[3]),
    .e(al_fff0fd72[0]),
    .o(al_e7bc5d6e));
  AL_MAP_LUT6 #(
    .EQN("(~F*(~(A)*(C*B)*~(D)*~(E)+A*(C*B)*~(D)*~(E)+~(A)*(C*B)*D*~(E)+A*(C*B)*D*~(E)+A*~((C*B))*~(D)*E+~(A)*(C*B)*~(D)*E+A*(C*B)*~(D)*E+A*~((C*B))*D*E+A*(C*B)*D*E))"),
    .INIT(64'h00000000aaeac0c0))
    al_2a3d05a (
    .a(al_e7bc5d6e),
    .b(al_32c99495[2]),
    .c(al_4e287126),
    .d(al_fff0fd72[0]),
    .e(al_fff0fd72[1]),
    .f(al_fff0fd72[2]),
    .o(al_471dc00c[0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_85dbf099 (
    .a(al_a21ad81c[0]),
    .b(al_a21ad81c[1]),
    .c(al_a21ad81c[2]),
    .d(al_a21ad81c[3]),
    .o(al_9ac9e635));
  AL_MAP_LUT6 #(
    .EQN("(~F*(~(A)*~((C*B))*D*~(E)+A*~((C*B))*D*~(E)+~(A)*~((C*B))*~(D)*E+A*~((C*B))*~(D)*E+~(A)*~((C*B))*D*E+~(A)*(C*B)*D*E))"),
    .INIT(64'h00000000553f3f00))
    al_217d02e6 (
    .a(al_9ac9e635),
    .b(al_32c99495[2]),
    .c(al_4e287126),
    .d(al_fff0fd72[0]),
    .e(al_fff0fd72[1]),
    .f(al_fff0fd72[2]),
    .o(al_471dc00c[1]));
  AL_MAP_LUT5 #(
    .EQN("(A*B*C*~(D)*~(E)+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E)"),
    .INIT(32'h03800080))
    al_3bbc8e7f (
    .a(al_9ac9e635),
    .b(al_fff0fd72[0]),
    .c(al_fff0fd72[1]),
    .d(al_fff0fd72[2]),
    .e(al_f6cc79fd),
    .o(al_471dc00c[2]));
  AL_DFF_X al_f0945f87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_acfeaf96[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_a21ad81c[0]));
  AL_DFF_X al_f971f9d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_acfeaf96[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_a21ad81c[1]));
  AL_DFF_X al_5c6c9496 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_acfeaf96[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_a21ad81c[2]));
  AL_DFF_X al_6ce2f8c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_acfeaf96[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_a21ad81c[3]));
  AL_DFF_X al_711f40b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_471dc00c[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_fff0fd72[0]));
  AL_DFF_X al_f9fcd693 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_471dc00c[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_fff0fd72[1]));
  AL_DFF_X al_5e875e6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_471dc00c[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_fff0fd72[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_cb87a87e (
    .a(al_7680352d),
    .b(al_278aa6ae[0]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[0]),
    .f(al_b05da9fd),
    .o(al_23bcf331[0]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_7ad4ea2a (
    .a(al_7680352d),
    .b(al_278aa6ae[10]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[10]),
    .f(al_b05da9fd),
    .o(al_23bcf331[10]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_42738fd6 (
    .a(al_7680352d),
    .b(al_278aa6ae[11]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[11]),
    .f(al_b05da9fd),
    .o(al_23bcf331[11]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_afde0ab0 (
    .a(al_278aa6ae[6]),
    .b(al_278aa6ae[7]),
    .c(al_278aa6ae[8]),
    .d(al_278aa6ae[9]),
    .e(al_278aa6ae[10]),
    .f(al_278aa6ae[11]),
    .o(al_17a2b8b));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_1a2242a2 (
    .a(al_278aa6ae[0]),
    .b(al_278aa6ae[1]),
    .c(al_278aa6ae[2]),
    .d(al_278aa6ae[3]),
    .e(al_278aa6ae[4]),
    .f(al_278aa6ae[5]),
    .o(al_da621072));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_aa4e0cd7 (
    .a(al_17a2b8b),
    .b(al_da621072),
    .c(al_278aa6ae[12]),
    .o(al_7680352d));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_d7a9769c (
    .a(al_7680352d),
    .b(al_278aa6ae[12]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[12]),
    .f(al_b05da9fd),
    .o(al_23bcf331[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_cf6232d5 (
    .a(al_7680352d),
    .b(al_278aa6ae[1]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[1]),
    .f(al_b05da9fd),
    .o(al_23bcf331[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_1a6a694e (
    .a(al_7680352d),
    .b(al_278aa6ae[2]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[2]),
    .f(al_b05da9fd),
    .o(al_23bcf331[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_97d4ab4c (
    .a(al_7680352d),
    .b(al_278aa6ae[3]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[3]),
    .f(al_b05da9fd),
    .o(al_23bcf331[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_a774e9d8 (
    .a(al_7680352d),
    .b(al_278aa6ae[4]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[4]),
    .f(al_b05da9fd),
    .o(al_23bcf331[4]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_1b8d157 (
    .a(al_7680352d),
    .b(al_278aa6ae[5]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[5]),
    .f(al_b05da9fd),
    .o(al_23bcf331[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_ee93a595 (
    .a(al_7680352d),
    .b(al_278aa6ae[6]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[6]),
    .f(al_b05da9fd),
    .o(al_23bcf331[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_e26b508f (
    .a(al_7680352d),
    .b(al_278aa6ae[7]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[7]),
    .f(al_b05da9fd),
    .o(al_23bcf331[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_9027ac29 (
    .a(al_7680352d),
    .b(al_278aa6ae[8]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[8]),
    .f(al_b05da9fd),
    .o(al_23bcf331[8]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~(D)*~(E)*~((~F*~A))+B*~(C)*~(D)*~(E)*~((~F*~A))+B*C*~(D)*~(E)*~((~F*~A))+B*~(C)*D*~(E)*~((~F*~A))+B*C*D*~(E)*~((~F*~A))+~(B)*~(C)*~(D)*E*~((~F*~A))+B*~(C)*~(D)*E*~((~F*~A))+B*C*~(D)*E*~((~F*~A))+B*~(C)*D*E*~((~F*~A))+B*C*D*E*~((~F*~A))+~(B)*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*~(D)*~(E)*(~F*~A)+B*~(C)*D*~(E)*(~F*~A)+B*C*D*~(E)*(~F*~A)+~(B)*~(C)*~(D)*E*(~F*~A)+B*~(C)*~(D)*E*(~F*~A)+~(B)*C*~(D)*E*(~F*~A)+B*C*~(D)*E*(~F*~A)+B*~(C)*D*E*(~F*~A)+B*C*D*E*(~F*~A))"),
    .INIT(64'hcccfcccfccdfcc8f))
    al_ba5e7c05 (
    .a(al_7680352d),
    .b(al_278aa6ae[9]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_56ef451f[9]),
    .f(al_b05da9fd),
    .o(al_23bcf331[9]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_4f239c8 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .o(al_c68f2ca9));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(~D*~B)))"),
    .INIT(16'ha0b0))
    al_5005247a (
    .a(al_ff9a0466),
    .b(al_278aa6ae[4]),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .o(al_3cb62398));
  AL_DFF_X al_8b5ddf4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3cb62398),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff9a0466));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_7c4281f0 (
    .a(al_73bb0740),
    .b(al_5e767b18),
    .c(al_5a579dd),
    .o(al_c5272fc1));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(32'h0000005c))
    al_b90e771a (
    .a(al_7680352d),
    .b(al_c5272fc1),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_b05da9fd),
    .o(al_fd60fee0[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*C*~(D)*~((~F*~E*B))+A*C*~(D)*(~F*~E*B)+~(A)*~(C)*D*(~F*~E*B)+A*~(C)*D*(~F*~E*B))"),
    .INIT(64'h00a000a000a00ca0))
    al_55bf95b3 (
    .a(al_7680352d),
    .b(al_73bb0740),
    .c(al_d2dd6034[0]),
    .d(al_d2dd6034[1]),
    .e(al_b05da9fd),
    .f(al_55ac2d11),
    .o(al_fd60fee0[1]));
  AL_DFF_X al_d098e861 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[8]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[8]));
  AL_DFF_X al_5510e75a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[9]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[9]));
  AL_DFF_X al_299723c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[10]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[10]));
  AL_DFF_X al_3b4bfabf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[11]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[11]));
  AL_DFF_X al_7a2dbcf2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[12]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[12]));
  AL_DFF_X al_8e18ad8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[0]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[0]));
  AL_DFF_X al_a7d3d2db (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[1]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[1]));
  AL_DFF_X al_141f0f0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[2]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[2]));
  AL_DFF_X al_3da2c8d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[3]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[3]));
  AL_DFF_X al_99f20154 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[4]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[4]));
  AL_DFF_X al_93dcfeeb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[5]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[5]));
  AL_DFF_X al_568e0bbc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[6]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[6]));
  AL_DFF_X al_501b56da (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_23bcf331[7]),
    .en(al_c68f2ca9),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_278aa6ae[7]));
  AL_DFF_X al_59b73838 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_fd60fee0[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d2dd6034[0]));
  AL_DFF_X al_14c602c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_fd60fee0[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d2dd6034[1]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_21d237d (
    .a(1'b0),
    .o({al_81a5ac08,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3cce3b84 (
    .a(al_278aa6ae[0]),
    .b(1'b1),
    .c(al_81a5ac08),
    .o({al_d424a202,al_56ef451f[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3ec977a8 (
    .a(al_278aa6ae[1]),
    .b(1'b0),
    .c(al_d424a202),
    .o({al_aaec830f,al_56ef451f[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_648c0a6f (
    .a(al_278aa6ae[2]),
    .b(1'b0),
    .c(al_aaec830f),
    .o({al_7680e48,al_56ef451f[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eb5e5000 (
    .a(al_278aa6ae[3]),
    .b(1'b0),
    .c(al_7680e48),
    .o({al_cb6844a5,al_56ef451f[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4a3926e3 (
    .a(al_278aa6ae[4]),
    .b(1'b0),
    .c(al_cb6844a5),
    .o({al_b53d4bb7,al_56ef451f[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6c223e2a (
    .a(al_278aa6ae[5]),
    .b(1'b0),
    .c(al_b53d4bb7),
    .o({al_1093568b,al_56ef451f[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1afe174f (
    .a(al_278aa6ae[6]),
    .b(1'b0),
    .c(al_1093568b),
    .o({al_720c32ab,al_56ef451f[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6378c461 (
    .a(al_278aa6ae[7]),
    .b(1'b0),
    .c(al_720c32ab),
    .o({al_cd4fb40c,al_56ef451f[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d761a780 (
    .a(al_278aa6ae[8]),
    .b(1'b0),
    .c(al_cd4fb40c),
    .o({al_174be6c3,al_56ef451f[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_de78356d (
    .a(al_278aa6ae[9]),
    .b(1'b0),
    .c(al_174be6c3),
    .o({al_24bcb54c,al_56ef451f[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a5c2f5ca (
    .a(al_278aa6ae[10]),
    .b(1'b0),
    .c(al_24bcb54c),
    .o({al_35d72057,al_56ef451f[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4c861fa6 (
    .a(al_278aa6ae[11]),
    .b(1'b0),
    .c(al_35d72057),
    .o({al_ef9c2399,al_56ef451f[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cca6dda1 (
    .a(al_278aa6ae[12]),
    .b(1'b0),
    .c(al_ef9c2399),
    .o({open_n11,al_56ef451f[12]}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_1b7bf60f (
    .a(al_c01774ad[0]),
    .b(al_7dd23876),
    .c(al_9c49a375[0]),
    .o(al_4228c99a[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_50b923ca (
    .a(al_c01774ad[1]),
    .b(al_7dd23876),
    .c(al_9c49a375[1]),
    .o(al_4228c99a[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_4b82007b (
    .a(al_c01774ad[2]),
    .b(al_7dd23876),
    .c(al_9c49a375[2]),
    .o(al_4228c99a[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_44fe290 (
    .a(al_c01774ad[3]),
    .b(al_7dd23876),
    .c(al_9c49a375[3]),
    .o(al_4228c99a[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_bb73e0e4 (
    .a(al_c01774ad[4]),
    .b(al_7dd23876),
    .c(al_9c49a375[4]),
    .o(al_4228c99a[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_a08a0302 (
    .a(al_c01774ad[5]),
    .b(al_7dd23876),
    .c(al_9c49a375[5]),
    .o(al_4228c99a[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_5f7b8a2b (
    .a(al_c01774ad[6]),
    .b(al_7dd23876),
    .c(al_9c49a375[6]),
    .o(al_4228c99a[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_15693db1 (
    .a(al_c01774ad[7]),
    .b(al_7dd23876),
    .c(al_9c49a375[7]),
    .o(al_4228c99a[7]));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_fdd14520 (
    .a(al_7dd23876),
    .b(al_32c99495[4]),
    .o(al_9ff01b51));
  AL_DFF_X al_95a29c0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9ff01b51),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_a231fc3f));
  AL_DFF_X al_7220ba86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(gmii_crs),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_4e287126));
  AL_DFF_X al_400d7df6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_32c99495[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_496839d3));
  AL_DFF_X al_e6eb8f1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_32c99495[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_5e767b18));
  AL_DFF_X al_9713360b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_32c99495[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_46f6a926));
  AL_DFF_X al_b052c3a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_32c99495[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1ea4ba5b));
  AL_DFF_X al_7c080a50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7b681f71),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_de9cd38));
  AL_DFF_X al_953d17cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b0d5abbb),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_b1d9ebd5));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~((~C*~B))*~(D)+A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*~((~C*~B))*D+~(A)*(~C*~B)*D)"),
    .INIT(16'h55fe))
    al_1a66e1a (
    .a(al_7fc110d7),
    .b(al_e11118e),
    .c(al_34e054a0),
    .d(al_c9168fb8[0]),
    .o(al_55a9d56d[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~((~C*~B))*~(D)*~(E)+A*~((~C*~B))*~(D)*~(E)+A*(~C*~B)*~(D)*~(E)+~(A)*~((~C*~B))*D*~(E)+~(A)*~((~C*~B))*~(D)*E+~(A)*(~C*~B)*~(D)*E+~(A)*~((~C*~B))*D*E+A*~((~C*~B))*D*E+~(A)*(~C*~B)*D*E+A*(~C*~B)*D*E)"),
    .INIT(32'hff5554fe))
    al_d9f7bf10 (
    .a(al_7fc110d7),
    .b(al_e11118e),
    .c(al_34e054a0),
    .d(al_c9168fb8[0]),
    .e(al_c9168fb8[1]),
    .o(al_55a9d56d[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~((~C*~B))*~((~E*~D))*~(F)+~(A)*~((~C*~B))*(~E*~D)*~(F)+A*~((~C*~B))*(~E*~D)*~(F)+A*(~C*~B)*(~E*~D)*~(F)+~(A)*~((~C*~B))*~((~E*~D))*F+A*~((~C*~B))*~((~E*~D))*F+~(A)*(~C*~B)*~((~E*~D))*F+A*(~C*~B)*~((~E*~D))*F+~(A)*~((~C*~B))*(~E*~D)*F+~(A)*(~C*~B)*(~E*~D)*F)"),
    .INIT(64'hffffff55545454fe))
    al_180839ef (
    .a(al_7fc110d7),
    .b(al_e11118e),
    .c(al_34e054a0),
    .d(al_c9168fb8[0]),
    .e(al_c9168fb8[1]),
    .f(al_c9168fb8[2]),
    .o(al_55a9d56d[2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~((~D*~C))*~(E)+A*~(B)*~((~D*~C))*~(E)+A*B*~((~D*~C))*~(E)+A*B*(~D*~C)*~(E)+~(A)*~(B)*~((~D*~C))*E+A*~(B)*~((~D*~C))*E+~(A)*B*~((~D*~C))*E+~(A)*~(B)*(~D*~C)*E+A*~(B)*(~D*~C)*E+~(A)*B*(~D*~C)*E)"),
    .INIT(32'h7777bbb8))
    al_ecfec970 (
    .a(al_f32db70e),
    .b(al_7fc110d7),
    .c(al_e11118e),
    .d(al_34e054a0),
    .e(al_c9168fb8[3]),
    .o(al_55a9d56d[3]));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~((~D*~C))*~((~E*A))*~(F)+~(B)*~((~D*~C))*(~E*A)*~(F)+B*~((~D*~C))*(~E*A)*~(F)+B*(~D*~C)*(~E*A)*~(F)+~(B)*~((~D*~C))*~((~E*A))*F+B*~((~D*~C))*~((~E*A))*F+~(B)*(~D*~C)*~((~E*A))*F+B*(~D*~C)*~((~E*A))*F+~(B)*~((~D*~C))*(~E*A)*F+~(B)*(~D*~C)*(~E*A)*F)"),
    .INIT(64'hffff77773330bbb8))
    al_590cd176 (
    .a(al_f32db70e),
    .b(al_7fc110d7),
    .c(al_e11118e),
    .d(al_34e054a0),
    .e(al_c9168fb8[3]),
    .f(al_c9168fb8[4]),
    .o(al_55a9d56d[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_c03c18dd (
    .a(al_7b30ef6a),
    .b(al_96ecb37f),
    .o(al_7fc110d7));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_2858e5af (
    .a(al_c9168fb8[0]),
    .b(al_c9168fb8[1]),
    .c(al_c9168fb8[2]),
    .o(al_f32db70e));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_6e121f6b (
    .a(al_f32db70e),
    .b(al_c9168fb8[3]),
    .c(al_c9168fb8[4]),
    .o(al_d4f4862c));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~((~D*~C))*~(E)+A*~(B)*~((~D*~C))*~(E)+A*B*~((~D*~C))*~(E)+A*B*(~D*~C)*~(E)+~(A)*~(B)*~((~D*~C))*E+A*~(B)*~((~D*~C))*E+~(A)*B*~((~D*~C))*E+~(A)*~(B)*(~D*~C)*E+A*~(B)*(~D*~C)*E+~(A)*B*(~D*~C)*E)"),
    .INIT(32'h7777bbb8))
    al_cb21f0fe (
    .a(al_d4f4862c),
    .b(al_7fc110d7),
    .c(al_e11118e),
    .d(al_34e054a0),
    .e(al_c9168fb8[5]),
    .o(al_55a9d56d[5]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_1607e503 (
    .a(al_c9168fb8[2]),
    .o(al_30c5253d[0]));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hf7b3))
    al_6ce5801e (
    .a(al_26eaf94a),
    .b(al_d7d3035f),
    .c(al_332a045d[0]),
    .d(al_cc156ef4[0]),
    .o(al_dbdaab6[0]));
  AL_MAP_LUT6 #(
    .EQN("~((B*A*~(E*D))*~(F)*~(C)+(B*A*~(E*D))*F*~(C)+~((B*A*~(E*D)))*F*C+(B*A*~(E*D))*F*C)"),
    .INIT(64'h0f070707fff7f7f7))
    al_1fb32657 (
    .a(al_aa981a62[4]),
    .b(al_5a579dd),
    .c(al_d7d3035f),
    .d(al_c9168fb8[4]),
    .e(al_c9168fb8[5]),
    .f(al_332a045d[10]),
    .o(al_537f614b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(C)*~((~D*B))*~(E)*~(F)+~(A)*C*~((~D*B))*~(E)*~(F)+~(A)*~(C)*(~D*B)*~(E)*~(F)+A*~(C)*(~D*B)*~(E)*~(F)+~(A)*C*(~D*B)*~(E)*~(F)+A*C*(~D*B)*~(E)*~(F)+~(A)*C*~((~D*B))*E*~(F)+~(A)*C*(~D*B)*E*~(F)+~(A)*~(C)*~((~D*B))*~(E)*F+~(A)*C*~((~D*B))*~(E)*F+~(A)*~(C)*(~D*B)*~(E)*F+A*~(C)*(~D*B)*~(E)*F+~(A)*C*(~D*B)*~(E)*F+A*C*(~D*B)*~(E)*F+~(A)*~(C)*~((~D*B))*E*F+A*~(C)*~((~D*B))*E*F+~(A)*C*~((~D*B))*E*F+~(A)*~(C)*(~D*B)*E*F+A*~(C)*(~D*B)*E*F+~(A)*C*(~D*B)*E*F)"),
    .INIT(64'h5f5f55dd505055dd))
    al_53414c5d (
    .a(al_537f614b),
    .b(al_ab37059b[1]),
    .c(al_26eaf94a),
    .d(al_5a579dd),
    .e(al_d7d3035f),
    .f(al_cc156ef4[10]),
    .o(al_dbdaab6[10]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    al_1bd29dec (
    .a(al_aa981a62[2]),
    .b(al_c9168fb8[3]),
    .c(al_c9168fb8[4]),
    .d(al_c9168fb8[5]),
    .o(al_ab37059b[2]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~(~D*~(C*B))))"),
    .INIT(32'h002aaaaa))
    al_82c56a11 (
    .a(al_aa981a62[5]),
    .b(al_c9168fb8[2]),
    .c(al_c9168fb8[3]),
    .d(al_c9168fb8[4]),
    .e(al_c9168fb8[5]),
    .o(al_ab37059b[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffacf0ac0fac00ac))
    al_7b54774c (
    .a(al_ab37059b[5]),
    .b(al_ab37059b[2]),
    .c(al_78564a3b),
    .d(al_d7d3035f),
    .e(al_332a045d[11]),
    .f(al_cc156ef4[11]),
    .o(al_dbdaab6[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_381fae22 (
    .a(al_ab37059b[3]),
    .b(al_ab37059b[6]),
    .c(al_5a579dd),
    .o(al_b06018b7));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hfa3aca0a))
    al_8d34b877 (
    .a(al_b06018b7),
    .b(al_26eaf94a),
    .c(al_d7d3035f),
    .d(al_332a045d[12]),
    .e(al_cc156ef4[12]),
    .o(al_dbdaab6[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    al_a2b54378 (
    .a(al_cf20ff1a),
    .b(al_aa981a62[7]),
    .c(al_c9168fb8[5]),
    .o(al_ab37059b[7]));
  AL_MAP_LUT6 #(
    .EQN("~((~B*A*~(E*D))*~(F)*~(C)+(~B*A*~(E*D))*F*~(C)+~((~B*A*~(E*D)))*F*C+(~B*A*~(E*D))*F*C)"),
    .INIT(64'h0f0d0d0dfffdfdfd))
    al_5981e7d7 (
    .a(al_aa981a62[4]),
    .b(al_5a579dd),
    .c(al_d7d3035f),
    .d(al_c9168fb8[4]),
    .e(al_c9168fb8[5]),
    .f(al_332a045d[13]),
    .o(al_f3a13de0));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~((D*A))*~(E)*~(F)+~(B)*C*~((D*A))*~(E)*~(F)+~(B)*~(C)*(D*A)*~(E)*~(F)+B*~(C)*(D*A)*~(E)*~(F)+~(B)*C*(D*A)*~(E)*~(F)+B*C*(D*A)*~(E)*~(F)+~(B)*C*~((D*A))*E*~(F)+~(B)*C*(D*A)*E*~(F)+~(B)*~(C)*~((D*A))*~(E)*F+~(B)*C*~((D*A))*~(E)*F+~(B)*~(C)*(D*A)*~(E)*F+B*~(C)*(D*A)*~(E)*F+~(B)*C*(D*A)*~(E)*F+B*C*(D*A)*~(E)*F+~(B)*~(C)*~((D*A))*E*F+B*~(C)*~((D*A))*E*F+~(B)*C*~((D*A))*E*F+~(B)*~(C)*(D*A)*E*F+B*~(C)*(D*A)*E*F+~(B)*C*(D*A)*E*F)"),
    .INIT(64'h3f3fbb333030bb33))
    al_4d9f9aef (
    .a(al_ab37059b[7]),
    .b(al_f3a13de0),
    .c(al_26eaf94a),
    .d(al_5a579dd),
    .e(al_d7d3035f),
    .f(al_cc156ef4[13]),
    .o(al_dbdaab6[13]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_dd74dbf4 (
    .a(al_aa981a62[8]),
    .b(al_c9168fb8[5]),
    .o(al_ab37059b[8]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffe2cce233e200e2))
    al_e5cb3b9d (
    .a(al_ab37059b[5]),
    .b(al_78564a3b),
    .c(al_ab37059b[8]),
    .d(al_d7d3035f),
    .e(al_332a045d[14]),
    .f(al_cc156ef4[14]),
    .o(al_dbdaab6[14]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_713889bf (
    .a(al_26eaf94a),
    .b(al_5a579dd),
    .c(al_d7d3035f),
    .o(al_78564a3b));
  AL_MAP_LUT5 #(
    .EQN("(~E*A*~(D*C*B))"),
    .INIT(32'h00002aaa))
    al_51dac1c3 (
    .a(al_aa981a62[9]),
    .b(al_c9168fb8[2]),
    .c(al_c9168fb8[3]),
    .d(al_c9168fb8[4]),
    .e(al_c9168fb8[5]),
    .o(al_ab37059b[9]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    al_d6938eb0 (
    .a(al_aa981a62[6]),
    .b(al_c9168fb8[3]),
    .c(al_c9168fb8[4]),
    .d(al_c9168fb8[5]),
    .o(al_ab37059b[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfafa0a0afc0cfc0c))
    al_1c9f0413 (
    .a(al_ab37059b[9]),
    .b(al_ab37059b[6]),
    .c(al_d7d3035f),
    .d(al_332a045d[15]),
    .e(al_cc156ef4[15]),
    .f(al_78564a3b),
    .o(al_dbdaab6[15]));
  AL_MAP_LUT6 #(
    .EQN("((~C*A)*~((F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B))*~(D)+(~C*A)*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*~(D)+~((~C*A))*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*D+(~C*A)*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*D)"),
    .INIT(64'hff0a330acc0a000a))
    al_f756f6e9 (
    .a(al_ab37059b[7]),
    .b(al_26eaf94a),
    .c(al_5a579dd),
    .d(al_d7d3035f),
    .e(al_332a045d[16]),
    .f(al_cc156ef4[16]),
    .o(al_dbdaab6[16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a4597b93 (
    .a(al_26eaf94a),
    .b(al_332a045d[17]),
    .c(al_cc156ef4[17]),
    .o(al_d991794b));
  AL_MAP_LUT5 #(
    .EQN("((~E*~C*B)*~(A)*~(D)+(~E*~C*B)*A*~(D)+~((~E*~C*B))*A*D+(~E*~C*B)*A*D)"),
    .INIT(32'haa00aa0c))
    al_cef3862 (
    .a(al_d991794b),
    .b(al_aa981a62[8]),
    .c(al_5a579dd),
    .d(al_d7d3035f),
    .e(al_c9168fb8[5]),
    .o(al_dbdaab6[17]));
  AL_MAP_LUT6 #(
    .EQN("((~C*A)*~((F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B))*~(D)+(~C*A)*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*~(D)+~((~C*A))*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*D+(~C*A)*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*D)"),
    .INIT(64'hff0a330acc0a000a))
    al_716051f5 (
    .a(al_ab37059b[9]),
    .b(al_26eaf94a),
    .c(al_5a579dd),
    .d(al_d7d3035f),
    .e(al_332a045d[18]),
    .f(al_cc156ef4[18]),
    .o(al_dbdaab6[18]));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hf7b3))
    al_f100fa9a (
    .a(al_26eaf94a),
    .b(al_d7d3035f),
    .c(al_332a045d[1]),
    .d(al_cc156ef4[1]),
    .o(al_dbdaab6[1]));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hf7b3))
    al_13ea8fb7 (
    .a(al_26eaf94a),
    .b(al_d7d3035f),
    .c(al_332a045d[2]),
    .d(al_cc156ef4[2]),
    .o(al_dbdaab6[2]));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hf7b3))
    al_b7096161 (
    .a(al_26eaf94a),
    .b(al_d7d3035f),
    .c(al_332a045d[3]),
    .d(al_cc156ef4[3]),
    .o(al_dbdaab6[3]));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hf7b3))
    al_a6105497 (
    .a(al_26eaf94a),
    .b(al_d7d3035f),
    .c(al_332a045d[4]),
    .d(al_cc156ef4[4]),
    .o(al_dbdaab6[4]));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hf7b3))
    al_fa10390a (
    .a(al_26eaf94a),
    .b(al_d7d3035f),
    .c(al_332a045d[5]),
    .d(al_cc156ef4[5]),
    .o(al_dbdaab6[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(C*~A)*~((F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B))*~(D)+~(C*~A)*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*~(D)+~(~(C*~A))*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*D+~(C*~A)*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*D)"),
    .INIT(64'hffaf33afccaf00af))
    al_44a8a3a2 (
    .a(al_aa981a62[0]),
    .b(al_26eaf94a),
    .c(al_5a579dd),
    .d(al_d7d3035f),
    .e(al_332a045d[6]),
    .f(al_cc156ef4[6]),
    .o(al_dbdaab6[6]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*D*C*B))"),
    .INIT(32'h2aaaaaaa))
    al_410ee15f (
    .a(al_aa981a62[1]),
    .b(al_c9168fb8[2]),
    .c(al_c9168fb8[3]),
    .d(al_c9168fb8[4]),
    .e(al_c9168fb8[5]),
    .o(al_ab37059b[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(C*~A)*~((F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B))*~(D)+~(C*~A)*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*~(D)+~(~(C*~A))*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*D+~(C*~A)*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*D)"),
    .INIT(64'hffaf33afccaf00af))
    al_e7fc111a (
    .a(al_ab37059b[1]),
    .b(al_26eaf94a),
    .c(al_5a579dd),
    .d(al_d7d3035f),
    .e(al_332a045d[7]),
    .f(al_cc156ef4[7]),
    .o(al_dbdaab6[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(C*~A)*~((F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B))*~(D)+~(C*~A)*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*~(D)+~(~(C*~A))*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*D+~(C*~A)*(F*~(E)*~(B)+F*E*~(B)+~(F)*E*B+F*E*B)*D)"),
    .INIT(64'hffaf33afccaf00af))
    al_9b97a414 (
    .a(al_ab37059b[2]),
    .b(al_26eaf94a),
    .c(al_5a579dd),
    .d(al_d7d3035f),
    .e(al_332a045d[8]),
    .f(al_cc156ef4[8]),
    .o(al_dbdaab6[8]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*D*~(~C*~B)))"),
    .INIT(32'h02aaaaaa))
    al_143ae0ce (
    .a(al_aa981a62[3]),
    .b(al_c9168fb8[2]),
    .c(al_c9168fb8[3]),
    .d(al_c9168fb8[4]),
    .e(al_c9168fb8[5]),
    .o(al_ab37059b[3]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfbf8cbc83b380b08))
    al_9385a1c0 (
    .a(al_ab37059b[3]),
    .b(al_78564a3b),
    .c(al_d7d3035f),
    .d(al_aa981a62[0]),
    .e(al_332a045d[9]),
    .f(al_cc156ef4[9]),
    .o(al_dbdaab6[9]));
  AL_DFF_X al_43e79bce (
    .ar(al_2dbca608),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ba6a9a7d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_26eaf94a));
  AL_MAP_LUT6 #(
    .EQN("(A*((~F*~E*~D)*~(B)*~(C)+(~F*~E*~D)*B*~(C)+~((~F*~E*~D))*B*C+(~F*~E*~D)*B*C))"),
    .INIT(64'h808080808080808a))
    al_c9bea1e8 (
    .a(al_143a100),
    .b(al_8ce032ae),
    .c(al_5a579dd),
    .d(al_332a045d[16]),
    .e(al_332a045d[17]),
    .f(al_332a045d[18]),
    .o(al_e7ec627));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    al_6bb02ac5 (
    .a(al_e7ec627),
    .b(tx_clk_en),
    .c(al_26eaf94a),
    .o(al_ba6a9a7d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_7e6d8384 (
    .a(al_332a045d[9]),
    .b(al_332a045d[10]),
    .c(al_332a045d[11]),
    .d(al_332a045d[12]),
    .e(al_332a045d[13]),
    .f(al_332a045d[14]),
    .o(al_459462b6));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_2ea9d888 (
    .a(al_459462b6),
    .b(tx_clk_en),
    .c(al_332a045d[0]),
    .d(al_332a045d[1]),
    .e(al_332a045d[3]),
    .f(al_332a045d[15]),
    .o(al_143a100));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_64921eaf (
    .a(al_332a045d[6]),
    .b(al_332a045d[7]),
    .c(al_332a045d[8]),
    .o(al_8ce032ae));
  AL_MAP_LUT4 #(
    .EQN("~(~D*A*~(~C*B))"),
    .INIT(16'hff5d))
    al_c0e40762 (
    .a(al_7521303d),
    .b(al_53f15a3f),
    .c(al_72f63008),
    .d(al_7b30ef6a),
    .o(al_ae71aa12));
  AL_DFF_X al_1e3b1811 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ae71aa12),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_53f15a3f));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_92a6176a (
    .a(al_26e8cb8e),
    .b(al_e29488b2[0]),
    .c(al_618d6d02[0]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_c05a6cac (
    .a(al_26e8cb8e),
    .b(al_e29488b2[10]),
    .c(al_618d6d02[10]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[10]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_ecdb0e06 (
    .a(al_26e8cb8e),
    .b(al_e29488b2[11]),
    .c(al_618d6d02[11]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[11]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_f13d191e (
    .a(al_26e8cb8e),
    .b(al_e29488b2[12]),
    .c(al_618d6d02[12]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[12]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_305ca31f (
    .a(al_26e8cb8e),
    .b(al_e29488b2[13]),
    .c(al_618d6d02[13]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[13]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_2882402a (
    .a(al_26e8cb8e),
    .b(al_e29488b2[1]),
    .c(al_618d6d02[1]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_4f2d3c83 (
    .a(al_26e8cb8e),
    .b(al_e29488b2[2]),
    .c(al_618d6d02[2]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[2]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_b2d32e3a (
    .a(al_26e8cb8e),
    .b(al_e29488b2[3]),
    .c(al_618d6d02[3]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_76324c75 (
    .a(al_26e8cb8e),
    .b(al_e29488b2[4]),
    .c(al_618d6d02[4]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_41d9f434 (
    .a(al_26e8cb8e),
    .b(al_e29488b2[5]),
    .c(al_618d6d02[5]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[5]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_f4f391ea (
    .a(al_26e8cb8e),
    .b(al_e29488b2[6]),
    .c(al_618d6d02[6]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[6]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_fee4efa3 (
    .a(al_26e8cb8e),
    .b(al_e29488b2[7]),
    .c(al_618d6d02[7]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_6a515646 (
    .a(al_26e8cb8e),
    .b(al_e29488b2[8]),
    .c(al_618d6d02[8]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[8]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    al_66a8ad47 (
    .a(al_26e8cb8e),
    .b(al_e29488b2[9]),
    .c(al_618d6d02[9]),
    .d(al_618d6d02[14]),
    .o(al_17c3d18e[9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_f43c5e0e (
    .a(al_1421d0c8),
    .b(al_ac2b4841),
    .c(al_7dd23876),
    .o(al_73bb0740));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_71865191 (
    .a(al_c9168fb8[2]),
    .b(al_c9168fb8[3]),
    .c(al_c9168fb8[4]),
    .o(al_cf20ff1a));
  AL_MAP_LUT6 #(
    .EQN("(E*B*~(C*~(~D*~(~F*A))))"),
    .INIT(64'h0ccc00000c4c0000))
    al_fdee4ebf (
    .a(al_cf20ff1a),
    .b(al_26eaf94a),
    .c(al_7b30ef6a),
    .d(al_ebd2d7),
    .e(al_d7d3035f),
    .f(al_c9168fb8[5]),
    .o(al_9ece8f02));
  AL_MAP_LUT6 #(
    .EQN("~(~(~F*D)*~(C*B*~(~E*~A)))"),
    .INIT(64'hc0c08080ffc0ff80))
    al_8e2a8b4b (
    .a(al_9ece8f02),
    .b(al_73bb0740),
    .c(al_496839d3),
    .d(al_3f0ffcfa),
    .e(al_e11118e),
    .f(al_618f3df7),
    .o(al_d42a4c18));
  AL_DFF_X al_3f35602 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d42a4c18),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3f0ffcfa));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_52f40e80 (
    .a(al_c8a3ac58),
    .b(al_7b30ef6a),
    .c(al_e9ae3746),
    .o(al_a8d42a04));
  AL_MAP_LUT6 #(
    .EQN("~(~(D*B)*~(F*~E*~(~C*A)))"),
    .INIT(64'hcc00fdf5cc00cc00))
    al_2b187a9 (
    .a(al_73bb0740),
    .b(al_a8d42a04),
    .c(al_adc2de29),
    .d(al_8c6e2d36),
    .e(al_6b8a9b19),
    .f(al_4024362),
    .o(al_3f77cd67));
  AL_DFF_X al_5a212df4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3f77cd67),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_8c6e2d36));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_d901acf2 (
    .a(al_c8a3ac58),
    .b(al_e9ae3746),
    .c(al_4024362),
    .o(al_f8ee3a1f));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_72db14b5 (
    .a(al_f8ee3a1f),
    .b(al_8c6e2d36),
    .c(al_266f6c4c),
    .d(al_2162c82e),
    .e(al_153acd6e),
    .o(al_3d1ba91a));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(~E*D)*~(~C*~B))"),
    .INIT(32'hababffab))
    al_90475776 (
    .a(al_bdf8d79f),
    .b(al_3d1ba91a),
    .c(al_73bb0740),
    .d(al_faa9857b),
    .e(al_618f3df7),
    .o(al_682de89f));
  AL_DFF_X al_769f2ee8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_682de89f),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_faa9857b));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(~D*~C*A))"),
    .INIT(16'hccce))
    al_c0f8eff9 (
    .a(al_f79b31c1),
    .b(al_266f6c4c),
    .c(al_e11118e),
    .d(al_618f3df7),
    .o(al_73642f31));
  AL_DFF_X al_b0ab5846 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_73642f31),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f79b31c1));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D*~B)*~(C*A))"),
    .INIT(32'hb3a0a0a0))
    al_a701968 (
    .a(al_a8d42a04),
    .b(al_8c6e2d36),
    .c(al_266f6c4c),
    .d(al_6b8a9b19),
    .e(al_4024362),
    .o(al_7b4de920));
  AL_DFF_X al_353eb613 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7b4de920),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_266f6c4c));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_ed7bdc74 (
    .a(al_f79b31c1),
    .b(al_6b8a9b19),
    .c(al_e9ae3746),
    .o(al_87c0c365));
  AL_DFF_X al_9efe00b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_87c0c365),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_b5c79ef6));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_2d103655 (
    .a(al_24ea5277),
    .b(al_eaafd789),
    .c(al_d567b233[0]),
    .o(al_e66356bf[0]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    al_8b3a13ad (
    .a(al_c98ce1a9),
    .b(al_eaafd789),
    .c(al_d62b96ee[2]),
    .o(al_e66356bf[10]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_8ce8bfd5 (
    .a(al_7b86230a),
    .b(al_d62b96ee[3]),
    .o(al_e66356bf[11]));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    al_2bde3d1e (
    .a(al_c560f884),
    .b(al_d567b233[5]),
    .c(al_d62b96ee[26]),
    .o(al_ebd48591));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*(C@B@A)))"),
    .INIT(32'h69ff9600))
    al_e52aa0d9 (
    .a(al_ebd48591),
    .b(al_24ea5277),
    .c(al_8f7895f1),
    .d(al_eaafd789),
    .e(al_d62b96ee[4]),
    .o(al_e66356bf[12]));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_67dc01ec (
    .a(al_d567b233[4]),
    .b(al_d567b233[5]),
    .c(al_d62b96ee[26]),
    .d(al_d62b96ee[27]),
    .o(al_c67dfcb5));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_b19f87a4 (
    .a(al_d567b233[1]),
    .b(al_d567b233[2]),
    .c(al_d62b96ee[29]),
    .d(al_d62b96ee[30]),
    .o(al_ac325ba1));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*(C@B@A)))"),
    .INIT(32'h69ff9600))
    al_500c90c3 (
    .a(al_c198e7cb),
    .b(al_c67dfcb5),
    .c(al_ac325ba1),
    .d(al_eaafd789),
    .e(al_d62b96ee[5]),
    .o(al_e66356bf[13]));
  AL_MAP_LUT6 #(
    .EQN("(E@(C*~(F@D@B@A)))"),
    .INIT(64'h6f9f90609f6f6090))
    al_402246b8 (
    .a(al_c67dfcb5),
    .b(al_2be5d117[0]),
    .c(al_eaafd789),
    .d(al_d567b233[3]),
    .e(al_d62b96ee[6]),
    .f(al_d62b96ee[28]),
    .o(al_e66356bf[14]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@E@D@C@A))"),
    .INIT(64'h8448488448848448))
    al_c9541b6 (
    .a(al_c560f884),
    .b(al_eaafd789),
    .c(al_d567b233[0]),
    .d(al_d567b233[4]),
    .e(al_d62b96ee[27]),
    .f(al_d62b96ee[31]),
    .o(al_8fda147c));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_f7c612fc (
    .a(al_8fda147c),
    .b(al_d62b96ee[7]),
    .o(al_e66356bf[15]));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(E@C@A)))"),
    .INIT(32'hb7487b84))
    al_60de22fb (
    .a(al_c560f884),
    .b(al_eaafd789),
    .c(al_d567b233[7]),
    .d(al_d62b96ee[8]),
    .e(al_d62b96ee[24]),
    .o(al_e66356bf[16]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_2ef5dfe2 (
    .a(al_ac325ba1),
    .b(al_8f7895f1),
    .c(al_eaafd789),
    .d(al_d62b96ee[9]),
    .o(al_e66356bf[17]));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(E@C@A)))"),
    .INIT(32'hb7487b84))
    al_9f33cdfa (
    .a(al_2be5d117[0]),
    .b(al_eaafd789),
    .c(al_d567b233[5]),
    .d(al_d62b96ee[10]),
    .e(al_d62b96ee[26]),
    .o(al_e66356bf[18]));
  AL_MAP_LUT6 #(
    .EQN("(D@(A*(F@E@C@B)))"),
    .INIT(64'hd7287d827d82d728))
    al_70afcf1d (
    .a(al_eaafd789),
    .b(al_d567b233[0]),
    .c(al_d567b233[4]),
    .d(al_d62b96ee[11]),
    .e(al_d62b96ee[27]),
    .f(al_d62b96ee[31]),
    .o(al_e66356bf[19]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_c5f3b56b (
    .a(al_bd399f0f),
    .b(al_eaafd789),
    .c(al_d567b233[1]),
    .o(al_e66356bf[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(D@B)))"),
    .INIT(16'h78d2))
    al_21be628a (
    .a(al_eaafd789),
    .b(al_d567b233[3]),
    .c(al_d62b96ee[12]),
    .d(al_d62b96ee[28]),
    .o(al_e66356bf[20]));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(D@B)))"),
    .INIT(16'h78d2))
    al_c1db0f77 (
    .a(al_eaafd789),
    .b(al_d567b233[2]),
    .c(al_d62b96ee[13]),
    .d(al_d62b96ee[29]),
    .o(al_e66356bf[21]));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(D@B)))"),
    .INIT(16'h78d2))
    al_bccbd3d2 (
    .a(al_eaafd789),
    .b(al_d567b233[7]),
    .c(al_d62b96ee[14]),
    .d(al_d62b96ee[24]),
    .o(al_e66356bf[22]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_32233c90 (
    .a(al_24ea5277),
    .b(al_8f7895f1),
    .c(al_eaafd789),
    .d(al_d62b96ee[15]),
    .o(al_e66356bf[23]));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(E@C@A)))"),
    .INIT(32'hb7487b84))
    al_2abc0c78 (
    .a(al_c198e7cb),
    .b(al_eaafd789),
    .c(al_d567b233[5]),
    .d(al_d62b96ee[16]),
    .e(al_d62b96ee[26]),
    .o(al_e66356bf[24]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    al_8282d0a4 (
    .a(al_c67dfcb5),
    .b(al_eaafd789),
    .c(al_d62b96ee[17]),
    .o(al_e66356bf[25]));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_9cbc5f7a (
    .a(al_d567b233[3]),
    .b(al_d567b233[4]),
    .c(al_d62b96ee[27]),
    .d(al_d62b96ee[28]),
    .o(al_abc33f01));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_6f8f9b52 (
    .a(al_24ea5277),
    .b(al_abc33f01),
    .c(al_eaafd789),
    .d(al_d62b96ee[18]),
    .o(al_e66356bf[26]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_3e3dc9bb (
    .a(al_c198e7cb),
    .b(al_c560f884),
    .c(al_eaafd789),
    .d(al_d62b96ee[19]),
    .o(al_e66356bf[27]));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(E@C@A)))"),
    .INIT(32'hb7487b84))
    al_10dbc41 (
    .a(al_ac325ba1),
    .b(al_eaafd789),
    .c(al_d567b233[5]),
    .d(al_d62b96ee[20]),
    .e(al_d62b96ee[26]),
    .o(al_e66356bf[28]));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(E@C@A)))"),
    .INIT(32'hb7487b84))
    al_ea2c75b0 (
    .a(al_2be5d117[0]),
    .b(al_eaafd789),
    .c(al_d567b233[4]),
    .d(al_d62b96ee[21]),
    .e(al_d62b96ee[27]),
    .o(al_e66356bf[29]));
  AL_MAP_LUT5 #(
    .EQN("(C*~((E@D@A))*~(B)+C*(E@D@A)*~(B)+~(C)*(E@D@A)*B+C*(E@D@A)*B)"),
    .INIT(32'hb87474b8))
    al_8ead4bd0 (
    .a(al_bd399f0f),
    .b(al_eaafd789),
    .c(al_d567b233[2]),
    .d(al_d567b233[5]),
    .e(al_d62b96ee[26]),
    .o(al_e66356bf[2]));
  AL_MAP_LUT6 #(
    .EQN("(D@(A*(F@E@C@B)))"),
    .INIT(64'hd7287d827d82d728))
    al_ab3effdb (
    .a(al_eaafd789),
    .b(al_d567b233[0]),
    .c(al_d567b233[3]),
    .d(al_d62b96ee[22]),
    .e(al_d62b96ee[28]),
    .f(al_d62b96ee[31]),
    .o(al_e66356bf[30]));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(D@B)))"),
    .INIT(16'h78d2))
    al_f9955ee1 (
    .a(al_eaafd789),
    .b(al_d567b233[2]),
    .c(al_d62b96ee[23]),
    .d(al_d62b96ee[29]),
    .o(al_e66356bf[31]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B@A))*~(C)+~D*(B@A)*~(C)+~(~D)*(B@A)*C+~D*(B@A)*C)"),
    .INIT(16'h9f90))
    al_e11da588 (
    .a(al_c198e7cb),
    .b(al_c67dfcb5),
    .c(al_eaafd789),
    .d(al_d567b233[3]),
    .o(al_e66356bf[3]));
  AL_MAP_LUT6 #(
    .EQN("(E*~((F@D@B@A))*~(C)+E*(F@D@B@A)*~(C)+~(E)*(F@D@B@A)*C+E*(F@D@B@A)*C)"),
    .INIT(64'h6f9f60909f6f9060))
    al_eeaa19ff (
    .a(al_24ea5277),
    .b(al_c67dfcb5),
    .c(al_eaafd789),
    .d(al_d567b233[3]),
    .e(al_d567b233[4]),
    .f(al_d62b96ee[28]),
    .o(al_e66356bf[4]));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_52df6da (
    .a(al_d567b233[1]),
    .b(al_d567b233[7]),
    .c(al_d62b96ee[24]),
    .d(al_d62b96ee[30]),
    .o(al_24ea5277));
  AL_MAP_LUT6 #(
    .EQN("(E*~((F@D@B@A))*~(C)+E*(F@D@B@A)*~(C)+~(E)*(F@D@B@A)*C+E*(F@D@B@A)*C)"),
    .INIT(64'h6f9f60909f6f9060))
    al_41d80115 (
    .a(al_bd399f0f),
    .b(al_c560f884),
    .c(al_eaafd789),
    .d(al_d567b233[4]),
    .e(al_d567b233[5]),
    .f(al_d62b96ee[27]),
    .o(al_e66356bf[5]));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_c4f37d14 (
    .a(al_d567b233[2]),
    .b(al_d567b233[3]),
    .c(al_d62b96ee[28]),
    .d(al_d62b96ee[29]),
    .o(al_c560f884));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_74c62764 (
    .a(al_d567b233[6]),
    .b(al_d62b96ee[25]),
    .o(al_8f7895f1));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    al_5e84ea72 (
    .a(al_8f7895f1),
    .b(al_d567b233[0]),
    .c(al_d62b96ee[31]),
    .o(al_c198e7cb));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_ff5bd3f0 (
    .a(al_c198e7cb),
    .b(al_24ea5277),
    .o(al_bd399f0f));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_492c0d98 (
    .a(al_d567b233[0]),
    .b(al_d567b233[1]),
    .c(al_d62b96ee[30]),
    .d(al_d62b96ee[31]),
    .o(al_2be5d117[0]));
  AL_MAP_LUT5 #(
    .EQN("(D@(C*~(E@B@A)))"),
    .INIT(32'h9f606f90))
    al_f9c990 (
    .a(al_ebd48591),
    .b(al_2be5d117[0]),
    .c(al_eaafd789),
    .d(al_d567b233[6]),
    .e(al_d62b96ee[25]),
    .o(al_e66356bf[6]));
  AL_MAP_LUT5 #(
    .EQN("(E@D@C@B@A)"),
    .INIT(32'h96696996))
    al_8b3e3aaf (
    .a(al_c67dfcb5),
    .b(al_d567b233[2]),
    .c(al_d567b233[7]),
    .d(al_d62b96ee[24]),
    .e(al_d62b96ee[29]),
    .o(al_c98ce1a9));
  AL_MAP_LUT5 #(
    .EQN("(D*~((E@C@A))*~(B)+D*(E@C@A)*~(B)+~(D)*(E@C@A)*B+D*(E@C@A)*B)"),
    .INIT(32'hb7847b48))
    al_c20e4d7e (
    .a(al_c98ce1a9),
    .b(al_eaafd789),
    .c(al_d567b233[0]),
    .d(al_d567b233[7]),
    .e(al_d62b96ee[31]),
    .o(al_e66356bf[7]));
  AL_MAP_LUT5 #(
    .EQN("(C*(E@D@B@A))"),
    .INIT(32'h60909060))
    al_12ef710b (
    .a(al_abc33f01),
    .b(al_8f7895f1),
    .c(al_eaafd789),
    .d(al_d567b233[7]),
    .e(al_d62b96ee[24]),
    .o(al_7b86230a));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_af47cfe8 (
    .a(al_7b86230a),
    .b(al_d62b96ee[0]),
    .o(al_e66356bf[8]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_ed97de70 (
    .a(al_ebd48591),
    .b(al_8f7895f1),
    .c(al_eaafd789),
    .d(al_d62b96ee[1]),
    .o(al_e66356bf[9]));
  AL_DFF_X al_5dd4b8e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[8]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[8]));
  AL_DFF_X al_cc174fe2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[9]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[9]));
  AL_DFF_X al_bfe3bc0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[10]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[10]));
  AL_DFF_X al_b7a791b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[11]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[11]));
  AL_DFF_X al_e17dab2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[12]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[12]));
  AL_DFF_X al_4f00245a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[13]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[13]));
  AL_DFF_X al_c80ea2e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[14]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[14]));
  AL_DFF_X al_c5095cf8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[15]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[15]));
  AL_DFF_X al_6da92d79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[16]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[16]));
  AL_DFF_X al_bc6b27e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[17]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[17]));
  AL_DFF_X al_823109e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[0]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[0]));
  AL_DFF_X al_bd16e50c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[18]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[18]));
  AL_DFF_X al_981eb9a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[19]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[19]));
  AL_DFF_X al_121a5065 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[20]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[20]));
  AL_DFF_X al_9afea46d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[21]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[21]));
  AL_DFF_X al_66977156 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[22]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[22]));
  AL_DFF_X al_239330dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[23]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[23]));
  AL_DFF_X al_24fd27e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[24]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[24]));
  AL_DFF_X al_d78bd415 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[25]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[25]));
  AL_DFF_X al_410ed77e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[26]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[26]));
  AL_DFF_X al_883a90bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[27]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[27]));
  AL_DFF_X al_4ab61b90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[1]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[1]));
  AL_DFF_X al_e261e5bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[28]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[28]));
  AL_DFF_X al_41909376 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[29]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[29]));
  AL_DFF_X al_9b8c495 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[30]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[30]));
  AL_DFF_X al_f4b5c3b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[31]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[31]));
  AL_DFF_X al_ad06e25a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[2]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[2]));
  AL_DFF_X al_b55b5cb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[3]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[3]));
  AL_DFF_X al_85f2d482 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[4]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[4]));
  AL_DFF_X al_3c5ece60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[5]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[5]));
  AL_DFF_X al_f6326f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[6]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[6]));
  AL_DFF_X al_c12f1cb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e66356bf[7]),
    .en(tx_clk_en),
    .sr(al_cb8cffb4[2]),
    .ss(1'b0),
    .q(al_d62b96ee[7]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_92042785 (
    .a(al_f5fd4d02),
    .b(al_931288d8[0]),
    .o(al_100aadd6));
  AL_DFF_X al_4ce79843 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_100aadd6),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eaafd789));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    al_85e5a1de (
    .a(al_c8a3ac58),
    .b(al_321109d3[0]),
    .o(al_aea1aa30[0]));
  AL_MAP_LUT3 #(
    .EQN("~(A*(C@B))"),
    .INIT(8'hd7))
    al_64c996bf (
    .a(al_c8a3ac58),
    .b(al_321109d3[0]),
    .c(al_321109d3[1]),
    .o(al_aea1aa30[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_58f10739 (
    .a(al_8c6e2d36),
    .b(al_c8a3ac58),
    .o(al_38320d7c));
  AL_DFF_X al_9124266f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_38320d7c),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9ba351db));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_56f4fe4 (
    .a(al_9953d0c8),
    .b(al_2ea27c82[1]),
    .o(al_d275691c[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_fe1b0c5f (
    .a(al_9953d0c8),
    .b(al_2ea27c82[3]),
    .o(al_d275691c[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_5f788706 (
    .a(al_9953d0c8),
    .b(al_2ea27c82[5]),
    .o(al_d275691c[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6f04371c (
    .a(al_9953d0c8),
    .b(al_1717406d),
    .c(al_2ea27c82[7]),
    .o(al_d275691c[7]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_dcff5cac (
    .a(al_9953d0c8),
    .b(al_2ea27c82[0]),
    .o(al_8b969422[0]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_6d13bfc6 (
    .a(al_9953d0c8),
    .b(al_2ea27c82[2]),
    .o(al_8b969422[2]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_323adb0a (
    .a(al_9953d0c8),
    .b(al_2ea27c82[4]),
    .o(al_8b969422[4]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_88ba83fa (
    .a(al_9953d0c8),
    .b(al_2ea27c82[6]),
    .o(al_8b969422[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A)*~((~C*~B))+D*A*~((~C*~B))+~(D)*A*(~C*~B)+D*A*(~C*~B))"),
    .INIT(16'hfe02))
    al_e63eebce (
    .a(al_3daf6177),
    .b(al_cd9f7a57),
    .c(al_bd8e6c56),
    .d(al_f5fe9553[0]),
    .o(al_da791a9b[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A)*~((~C*~B))+D*A*~((~C*~B))+~(D)*A*(~C*~B)+D*A*(~C*~B))"),
    .INIT(16'hfe02))
    al_c0c531c8 (
    .a(al_3daf6177),
    .b(al_cd9f7a57),
    .c(al_bd8e6c56),
    .d(al_f5fe9553[1]),
    .o(al_da791a9b[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A)*~((~C*~B))+D*A*~((~C*~B))+~(D)*A*(~C*~B)+D*A*(~C*~B))"),
    .INIT(16'hfe02))
    al_ff1db8ff (
    .a(al_3daf6177),
    .b(al_cd9f7a57),
    .c(al_bd8e6c56),
    .d(al_f5fe9553[2]),
    .o(al_da791a9b[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A)*~((~C*~B))+D*A*~((~C*~B))+~(D)*A*(~C*~B)+D*A*(~C*~B))"),
    .INIT(16'hfe02))
    al_85f8a93 (
    .a(al_3daf6177),
    .b(al_cd9f7a57),
    .c(al_bd8e6c56),
    .d(al_f5fe9553[3]),
    .o(al_da791a9b[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_683a52fc (
    .a(al_cd9f7a57),
    .b(al_bd8e6c56),
    .c(al_f5fe9553[4]),
    .o(al_da791a9b[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_bec6f123 (
    .a(al_cd9f7a57),
    .b(al_bd8e6c56),
    .c(al_f5fe9553[5]),
    .o(al_da791a9b[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_d6114269 (
    .a(al_cd9f7a57),
    .b(al_bd8e6c56),
    .c(al_f5fe9553[6]),
    .o(al_da791a9b[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_b39024f3 (
    .a(al_cd9f7a57),
    .b(al_bd8e6c56),
    .c(al_f5fe9553[7]),
    .o(al_da791a9b[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d5f772bd (
    .a(al_f5fd4d02),
    .b(al_31841a5b[0]),
    .o(al_47ab7609[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_4c52647b (
    .a(al_f5fd4d02),
    .b(al_31841a5b[1]),
    .o(al_47ab7609[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_aa8910b4 (
    .a(al_f5fd4d02),
    .b(al_31841a5b[2]),
    .o(al_47ab7609[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d4736001 (
    .a(al_f5fd4d02),
    .b(al_31841a5b[3]),
    .o(al_47ab7609[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_7be9026b (
    .a(al_f5fd4d02),
    .b(al_31841a5b[4]),
    .o(al_47ab7609[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f6592672 (
    .a(al_f5fd4d02),
    .b(al_31841a5b[5]),
    .o(al_47ab7609[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f3654e4e (
    .a(al_f5fd4d02),
    .b(al_31841a5b[6]),
    .o(al_47ab7609[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_696447d3 (
    .a(al_f5fd4d02),
    .b(al_31841a5b[7]),
    .o(al_47ab7609[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_a7f2283c (
    .a(al_7b30ef6a),
    .b(al_d567b233[0]),
    .o(al_d1fcb50b[0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .INIT(16'hfe32))
    al_fccc7769 (
    .a(al_d1fcb50b[0]),
    .b(al_9ba351db),
    .c(al_3daf6177),
    .d(al_d62b96ee[31]),
    .o(al_f24f9b58[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_8d9eaf5a (
    .a(al_7b30ef6a),
    .b(al_d567b233[1]),
    .o(al_d1fcb50b[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .INIT(16'hfe32))
    al_cdf2c29b (
    .a(al_d1fcb50b[1]),
    .b(al_9ba351db),
    .c(al_3daf6177),
    .d(al_d62b96ee[30]),
    .o(al_f24f9b58[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b0559368 (
    .a(al_7b30ef6a),
    .b(al_d567b233[2]),
    .o(al_d1fcb50b[2]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .INIT(16'hfe32))
    al_aa8212cf (
    .a(al_d1fcb50b[2]),
    .b(al_9ba351db),
    .c(al_3daf6177),
    .d(al_d62b96ee[29]),
    .o(al_f24f9b58[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_fed4c718 (
    .a(al_7b30ef6a),
    .b(al_d567b233[3]),
    .o(al_d1fcb50b[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .INIT(16'hfe32))
    al_456e5ad7 (
    .a(al_d1fcb50b[3]),
    .b(al_9ba351db),
    .c(al_3daf6177),
    .d(al_d62b96ee[28]),
    .o(al_f24f9b58[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_3c4dd286 (
    .a(al_7b30ef6a),
    .b(al_d567b233[4]),
    .o(al_d1fcb50b[4]));
  AL_MAP_LUT4 #(
    .EQN("((~C*A)*~(D)*~(B)+(~C*A)*D*~(B)+~((~C*A))*D*B+(~C*A)*D*B)"),
    .INIT(16'hce02))
    al_e418dd6 (
    .a(al_d1fcb50b[4]),
    .b(al_9ba351db),
    .c(al_3daf6177),
    .d(al_d62b96ee[27]),
    .o(al_f24f9b58[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c6993a89 (
    .a(al_7b30ef6a),
    .b(al_d567b233[5]),
    .o(al_d1fcb50b[5]));
  AL_MAP_LUT4 #(
    .EQN("((~C*A)*~(D)*~(B)+(~C*A)*D*~(B)+~((~C*A))*D*B+(~C*A)*D*B)"),
    .INIT(16'hce02))
    al_d4621067 (
    .a(al_d1fcb50b[5]),
    .b(al_9ba351db),
    .c(al_3daf6177),
    .d(al_d62b96ee[26]),
    .o(al_f24f9b58[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_dca910ec (
    .a(al_7b30ef6a),
    .b(al_d567b233[6]),
    .o(al_d1fcb50b[6]));
  AL_MAP_LUT4 #(
    .EQN("((~C*A)*~(D)*~(B)+(~C*A)*D*~(B)+~((~C*A))*D*B+(~C*A)*D*B)"),
    .INIT(16'hce02))
    al_60c687f9 (
    .a(al_d1fcb50b[6]),
    .b(al_9ba351db),
    .c(al_3daf6177),
    .d(al_d62b96ee[25]),
    .o(al_f24f9b58[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_1d5f08e1 (
    .a(al_7b30ef6a),
    .b(al_d567b233[7]),
    .o(al_d1fcb50b[7]));
  AL_MAP_LUT4 #(
    .EQN("((~C*A)*~(D)*~(B)+(~C*A)*D*~(B)+~((~C*A))*D*B+(~C*A)*D*B)"),
    .INIT(16'hce02))
    al_a6df5d9b (
    .a(al_d1fcb50b[7]),
    .b(al_9ba351db),
    .c(al_3daf6177),
    .d(al_d62b96ee[24]),
    .o(al_f24f9b58[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_829d8c0a (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[0]),
    .o(al_49200bab[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_8596e244 (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[10]),
    .o(al_49200bab[10]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_9820fbaf (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[11]),
    .o(al_49200bab[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_b541bc47 (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[12]),
    .o(al_49200bab[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_14acd619 (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[13]),
    .o(al_49200bab[13]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h8f07))
    al_5e89a1aa (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_5a579dd),
    .d(al_83a6bf62[14]),
    .o(al_49200bab[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_7888136f (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[1]),
    .o(al_49200bab[1]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_b1ffd33a (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[2]),
    .o(al_49200bab[2]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h8f07))
    al_b533933f (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_5a579dd),
    .d(al_83a6bf62[3]),
    .o(al_49200bab[3]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D)*~((B*A))+C*D*~((B*A))+~(C)*D*(B*A)+C*D*(B*A))"),
    .INIT(16'hf870))
    al_f601eb25 (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_5a579dd),
    .d(al_83a6bf62[4]),
    .o(al_49200bab[4]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    .INIT(16'h8f07))
    al_2a687a91 (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_5a579dd),
    .d(al_83a6bf62[5]),
    .o(al_49200bab[5]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_147ab3ae (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[6]),
    .o(al_49200bab[6]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_d0e86122 (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[7]),
    .o(al_49200bab[7]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_49ee0e0d (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[8]),
    .o(al_49200bab[8]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_ec7361d6 (
    .a(al_3f0ffcfa),
    .b(al_cd3c4af6),
    .c(al_83a6bf62[9]),
    .o(al_49200bab[9]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_aa21cd92 (
    .a(al_3f0ffcfa),
    .b(al_e11118e),
    .c(al_618f3df7),
    .o(al_9ce6a803));
  AL_DFF_X al_d6165720 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9ce6a803),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f6cc79fd));
  AL_DFF_X al_4e6b1d27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d8e2b166),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4bdde34));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_5c3fb935 (
    .a(al_2453f186[1]),
    .b(al_2453f186[2]),
    .c(al_2453f186[3]),
    .d(al_2453f186[4]),
    .e(al_2453f186[5]),
    .f(al_2453f186[6]),
    .o(al_f2be847d));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_6009b8a2 (
    .a(al_f2be847d),
    .b(al_6f12ed1d),
    .c(al_2453f186[0]),
    .d(al_2453f186[7]),
    .o(al_6becface));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(A)*~((E*B))+D*A*~((E*B))+~(D)*A*(E*B)+D*A*(E*B)))"),
    .INIT(32'h0b080f00))
    al_55be8f99 (
    .a(al_6becface),
    .b(tx_clk_en),
    .c(al_2dbca608),
    .d(al_4bdde34),
    .e(al_cb8cffb4[4]),
    .o(al_d8e2b166));
  AL_DFF_X al_5975185b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8eaf8008),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_136addab));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_17d1ca35 (
    .a(al_d567b233[1]),
    .b(al_d567b233[2]),
    .c(al_d567b233[3]),
    .d(al_d567b233[4]),
    .e(al_d567b233[5]),
    .f(al_d567b233[6]),
    .o(al_22412e0c));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_d3332f80 (
    .a(al_22412e0c),
    .b(al_6f12ed1d),
    .c(al_d567b233[0]),
    .d(al_d567b233[7]),
    .o(al_c2479eab));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(A)*~((E*B))+D*A*~((E*B))+~(D)*A*(E*B)+D*A*(E*B)))"),
    .INIT(32'h0b080f00))
    al_8e4b4f24 (
    .a(al_c2479eab),
    .b(tx_clk_en),
    .c(al_2dbca608),
    .d(al_136addab),
    .e(al_cb8cffb4[4]),
    .o(al_8eaf8008));
  AL_DFF_X al_b5338440 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4210af67),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9c0fa32));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_f9d49d0e (
    .a(al_31841a5b[1]),
    .b(al_31841a5b[2]),
    .c(al_31841a5b[3]),
    .d(al_31841a5b[4]),
    .e(al_31841a5b[5]),
    .f(al_31841a5b[6]),
    .o(al_2be5cde7));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_fcf7593a (
    .a(al_2be5cde7),
    .b(al_6f12ed1d),
    .c(al_31841a5b[0]),
    .d(al_31841a5b[7]),
    .o(al_c2428aac));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(A)*~((E*B))+D*A*~((E*B))+~(D)*A*(E*B)+D*A*(E*B)))"),
    .INIT(32'h0b080f00))
    al_9ae811b0 (
    .a(al_c2428aac),
    .b(tx_clk_en),
    .c(al_2dbca608),
    .d(al_c9c0fa32),
    .e(al_cb8cffb4[4]),
    .o(al_4210af67));
  AL_DFF_X al_e80260fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_279abee0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8e6107a7));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_c33e9668 (
    .a(al_f5fe9553[1]),
    .b(al_f5fe9553[2]),
    .c(al_f5fe9553[3]),
    .d(al_f5fe9553[4]),
    .e(al_f5fe9553[5]),
    .f(al_f5fe9553[6]),
    .o(al_b8bd8e77));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_e00f3578 (
    .a(al_b8bd8e77),
    .b(al_6f12ed1d),
    .c(al_f5fe9553[0]),
    .d(al_f5fe9553[7]),
    .o(al_32c6ecc7));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(A)*~((E*B))+D*A*~((E*B))+~(D)*A*(E*B)+D*A*(E*B)))"),
    .INIT(32'h0b080f00))
    al_c8b53959 (
    .a(al_32c6ecc7),
    .b(tx_clk_en),
    .c(al_2dbca608),
    .d(al_8e6107a7),
    .e(al_cb8cffb4[4]),
    .o(al_279abee0));
  AL_DFF_X al_de3af54e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f78cc6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15bf91ee));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(A)*~((E*B))+D*A*~((E*B))+~(D)*A*(E*B)+D*A*(E*B)))"),
    .INIT(32'h0b080f00))
    al_baa77f8e (
    .a(al_d73f3ba1),
    .b(tx_clk_en),
    .c(al_2dbca608),
    .d(al_15bf91ee),
    .e(al_cb8cffb4[4]),
    .o(al_1f78cc6));
  AL_DFF_X al_7c24ce29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b42ee6d4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af4842d7));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_7318be50 (
    .a(al_2ea27c82[1]),
    .b(al_2ea27c82[2]),
    .c(al_2ea27c82[3]),
    .d(al_2ea27c82[4]),
    .e(al_2ea27c82[5]),
    .f(al_2ea27c82[6]),
    .o(al_856accff));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_878bebee (
    .a(al_856accff),
    .b(al_6f12ed1d),
    .c(al_2ea27c82[0]),
    .d(al_2ea27c82[7]),
    .o(al_d73f3ba1));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(A)*~((E*B))+D*A*~((E*B))+~(D)*A*(E*B)+D*A*(E*B)))"),
    .INIT(32'h0b080f00))
    al_a6068e49 (
    .a(al_d73f3ba1),
    .b(tx_clk_en),
    .c(al_2dbca608),
    .d(al_af4842d7),
    .e(al_cb8cffb4[5]),
    .o(al_b42ee6d4));
  AL_DFF_X al_8c4012f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4952d975),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_336bd542));
  AL_MAP_LUT5 #(
    .EQN("(~B*(C*~(E)*~((D*A))+C*E*~((D*A))+~(C)*E*(D*A)+C*E*(D*A)))"),
    .INIT(32'h32301030))
    al_439ec926 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_336bd542),
    .d(al_cb8cffb4[4]),
    .e(al_2453f186[0]),
    .o(al_4952d975));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D@(~B*~A)))"),
    .INIT(16'h10e0))
    al_4f9f5bc4 (
    .a(al_3fc75a33),
    .b(al_b241735d),
    .c(al_8a331b5c),
    .d(al_1b8c3389[0]),
    .o(al_ee979a13[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_ca411be (
    .a(al_1b8c3389[0]),
    .b(al_1b8c3389[1]),
    .c(al_1b8c3389[2]),
    .d(al_1b8c3389[3]),
    .o(al_c75b827e));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~(C*~B*~A))"),
    .INIT(32'hef000000))
    al_d9adfc09 (
    .a(al_e5994b5e),
    .b(al_b241735d),
    .c(al_a2667927),
    .d(al_c75b827e),
    .e(al_1b8c3389[4]),
    .o(al_c89ba6ec));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_67511136 (
    .a(al_1b8c3389[5]),
    .b(al_1b8c3389[6]),
    .c(al_1b8c3389[7]),
    .d(al_1b8c3389[8]),
    .o(al_19aaf769));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_a7aad90f (
    .a(al_c89ba6ec),
    .b(al_8a331b5c),
    .c(al_19aaf769),
    .d(al_1b8c3389[9]),
    .e(al_1b8c3389[10]),
    .o(al_ee979a13[10]));
  AL_MAP_LUT5 #(
    .EQN("(C*(E@(D*~(~B*~A))))"),
    .INIT(32'h10f0e000))
    al_239e5cee (
    .a(al_3fc75a33),
    .b(al_b241735d),
    .c(al_8a331b5c),
    .d(al_1b8c3389[0]),
    .e(al_1b8c3389[1]),
    .o(al_ee979a13[1]));
  AL_MAP_LUT6 #(
    .EQN("(C*(F@(E*D*~(~B*~A))))"),
    .INIT(64'h10f0f0f0e0000000))
    al_2740e85e (
    .a(al_3fc75a33),
    .b(al_b241735d),
    .c(al_8a331b5c),
    .d(al_1b8c3389[0]),
    .e(al_1b8c3389[1]),
    .f(al_1b8c3389[2]),
    .o(al_ee979a13[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_e0c82066 (
    .a(al_1b8c3389[0]),
    .b(al_1b8c3389[1]),
    .c(al_1b8c3389[2]),
    .o(al_3009e595));
  AL_MAP_LUT5 #(
    .EQN("(C*(E@(D*~(~B*~A))))"),
    .INIT(32'h10f0e000))
    al_5705394d (
    .a(al_3fc75a33),
    .b(al_b241735d),
    .c(al_8a331b5c),
    .d(al_3009e595),
    .e(al_1b8c3389[3]),
    .o(al_ee979a13[3]));
  AL_MAP_LUT5 #(
    .EQN("(C*(E@(D*~(~B*~A))))"),
    .INIT(32'h10f0e000))
    al_977df0c5 (
    .a(al_3fc75a33),
    .b(al_b241735d),
    .c(al_8a331b5c),
    .d(al_c75b827e),
    .e(al_1b8c3389[4]),
    .o(al_ee979a13[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_fc62c6fe (
    .a(al_c89ba6ec),
    .b(al_8a331b5c),
    .c(al_1b8c3389[5]),
    .o(al_ee979a13[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_d0a2cf52 (
    .a(al_c89ba6ec),
    .b(al_8a331b5c),
    .c(al_1b8c3389[5]),
    .d(al_1b8c3389[6]),
    .o(al_ee979a13[6]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_6e5faf4 (
    .a(al_c89ba6ec),
    .b(al_8a331b5c),
    .c(al_1b8c3389[5]),
    .d(al_1b8c3389[6]),
    .e(al_1b8c3389[7]),
    .o(al_ee979a13[7]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@(E*D*C*A)))"),
    .INIT(64'h4ccccccc80000000))
    al_c771a619 (
    .a(al_c89ba6ec),
    .b(al_8a331b5c),
    .c(al_1b8c3389[5]),
    .d(al_1b8c3389[6]),
    .e(al_1b8c3389[7]),
    .f(al_1b8c3389[8]),
    .o(al_ee979a13[8]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_77a1c58c (
    .a(al_c89ba6ec),
    .b(al_8a331b5c),
    .c(al_19aaf769),
    .d(al_1b8c3389[9]),
    .o(al_ee979a13[9]));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*A)"),
    .INIT(32'h20000000))
    al_62166d47 (
    .a(al_7521303d),
    .b(al_53f15a3f),
    .c(al_846b6533),
    .d(al_6f12ed1d),
    .e(al_b4f442b4),
    .o(al_adae5a89));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_188ee755 (
    .a(al_e11118e),
    .b(al_cd9f7a57),
    .c(al_49948f6),
    .d(al_d7d3035f),
    .o(al_a51573d2));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~C*~A*~(E*D)))"),
    .INIT(32'hccc8c8c8))
    al_aaa841f7 (
    .a(al_adae5a89),
    .b(al_a51573d2),
    .c(al_72f63008),
    .d(al_7694b99f),
    .e(al_24faf4d6),
    .o(al_5563a8fd));
  AL_DFF_X al_529e89bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5563a8fd),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_72f63008));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*~A)"),
    .INIT(64'h0000000000000004))
    al_b09c804f (
    .a(al_72f63008),
    .b(al_846b6533),
    .c(al_7694b99f),
    .d(al_e11118e),
    .e(al_153acd6e),
    .f(al_49948f6),
    .o(al_77e56b3a));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~((C*~B))*~(D)*~(E)+~(A)*~((C*~B))*D*~(E)+~(A)*~((C*~B))*~(D)*E+A*~((C*~B))*~(D)*E+~(A)*~((C*~B))*D*E+A*~((C*~B))*D*E+~(A)*(C*~B)*D*E+A*(C*~B)*D*E)"),
    .INIT(32'hffcf4545))
    al_1b28facc (
    .a(al_53f15a3f),
    .b(al_f79b31c1),
    .c(al_6f12ed1d),
    .d(al_2162c82e),
    .e(al_24faf4d6),
    .o(al_807f5a12));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*C*~B)*~(~E*A))"),
    .INIT(32'h3000baaa))
    al_ff9f79da (
    .a(al_77e56b3a),
    .b(al_807f5a12),
    .c(al_7521303d),
    .d(al_e9ae3746),
    .e(al_d7d3035f),
    .o(al_9a1b441a));
  AL_DFF_X al_272ed2e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9a1b441a),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_846b6533));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    al_ab99f057 (
    .a(al_72f63008),
    .b(al_7694b99f),
    .c(al_49948f6),
    .d(al_d7d3035f),
    .o(al_67f58f23));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    al_86690d3e (
    .a(al_67f58f23),
    .b(al_7521303d),
    .c(al_53f15a3f),
    .d(al_846b6533),
    .e(al_b4f442b4),
    .o(al_3deafd60));
  AL_DFF_X al_97618564 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3deafd60),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_7694b99f));
  AL_MAP_LUT6 #(
    .EQN("(C*~(~F*~E)*~(~B*~(D*A)))"),
    .INIT(64'he0c0e0c0e0c00000))
    al_c663ccd2 (
    .a(al_8c6e2d36),
    .b(al_266f6c4c),
    .c(al_803bd5d9),
    .d(al_b96742e9),
    .e(al_321109d3[0]),
    .f(al_321109d3[1]),
    .o(al_4ab17dc7));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(~D*B)))"),
    .INIT(16'h0a0e))
    al_797c0941 (
    .a(al_4ab17dc7),
    .b(al_c8a3ac58),
    .c(al_7b30ef6a),
    .d(al_e9ae3746),
    .o(al_46a6aa32));
  AL_DFF_X al_2520d759 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_46a6aa32),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c8a3ac58));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_1f4331d6 (
    .a(al_c8a3ac58),
    .b(al_321109d3[0]),
    .c(al_321109d3[1]),
    .o(al_376757cc));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*B*A))"),
    .INIT(16'h070f))
    al_a0e88213 (
    .a(al_376757cc),
    .b(al_f79b31c1),
    .c(al_f718b05a),
    .d(al_6b8a9b19),
    .o(al_83146215));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(B*~A*~(~D*C)))"),
    .INIT(32'h0000bbfb))
    al_dce97d5 (
    .a(al_bdf8d79f),
    .b(al_83146215),
    .c(al_266f6c4c),
    .d(al_803bd5d9),
    .e(al_153acd6e),
    .o(al_53f06a44));
  AL_DFF_X al_67757230 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_53f06a44),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f718b05a));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_503a99b8 (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[0]),
    .c(al_5305cb61[0]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_e907d01f (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[10]),
    .c(al_5305cb61[10]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[10]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_cc50479a (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[11]),
    .c(al_5305cb61[11]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[11]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_c23bde93 (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[12]),
    .c(al_5305cb61[12]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[12]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_124a34c9 (
    .a(al_8c6e2d36),
    .b(al_846b6533),
    .c(al_7694b99f),
    .d(al_c8a3ac58),
    .e(al_4024362),
    .o(al_c710cf1a));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_1c83d228 (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[13]),
    .c(al_5305cb61[13]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[13]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    al_e172e7e4 (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[14]),
    .c(al_5305cb61[14]),
    .o(al_b084da19[14]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_9e191dcf (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[1]),
    .c(al_5305cb61[1]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[1]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(E)+C*D*~(E)+~(C)*D*E+C*D*E)*~(B)*~(A)+(C*~(D)*~(E)+C*D*~(E)+~(C)*D*E+C*D*E)*B*~(A)+~((C*~(D)*~(E)+C*D*~(E)+~(C)*D*E+C*D*E))*B*A+(C*~(D)*~(E)+C*D*~(E)+~(C)*D*E+C*D*E)*B*A)"),
    .INIT(32'hdd88d8d8))
    al_abe66acc (
    .a(al_c710cf1a),
    .b(al_803bd5d9),
    .c(al_b7d1cff2[2]),
    .d(al_5305cb61[2]),
    .e(al_5305cb61[14]),
    .o(al_b084da19[2]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_d54783df (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[3]),
    .c(al_5305cb61[3]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[3]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_32235768 (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[4]),
    .c(al_5305cb61[4]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[4]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_34ab977 (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[5]),
    .c(al_5305cb61[5]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[5]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_275f0979 (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[6]),
    .c(al_5305cb61[6]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[6]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_3abd5f1a (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[7]),
    .c(al_5305cb61[7]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[7]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_e174f006 (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[8]),
    .c(al_5305cb61[8]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[8]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    al_fc3bb1cf (
    .a(al_c710cf1a),
    .b(al_b7d1cff2[9]),
    .c(al_5305cb61[9]),
    .d(al_5305cb61[14]),
    .o(al_b084da19[9]));
  AL_MAP_LUT6 #(
    .EQN("~((F*B)*~((A*~(E*C)))*~(D)+(F*B)*(A*~(E*C))*~(D)+~((F*B))*(A*~(E*C))*D+(F*B)*(A*~(E*C))*D)"),
    .INIT(64'hf5335533f5ff55ff))
    al_c5645713 (
    .a(al_376757cc),
    .b(al_8c6e2d36),
    .c(al_f79b31c1),
    .d(al_803bd5d9),
    .e(al_6b8a9b19),
    .f(al_b96742e9),
    .o(al_cf358e1e));
  AL_MAP_LUT6 #(
    .EQN("~(A*~(~F*~E*D*~C*~B))"),
    .INIT(64'h5555555555555755))
    al_8055c045 (
    .a(al_cf358e1e),
    .b(al_72f63008),
    .c(al_7694b99f),
    .d(al_3d294c28),
    .e(al_7b30ef6a),
    .f(al_153acd6e),
    .o(al_a5c6fbcc));
  AL_DFF_X al_b23c98ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a5c6fbcc),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3d294c28));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_b921583a (
    .a(al_73bb0740),
    .b(al_7521303d),
    .o(al_e5bd99ae));
  AL_DFF_X al_6d84b16e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e5bd99ae),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9aa134ca));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_d88b66c8 (
    .a(al_eb2b30c3[8]),
    .b(al_eb2b30c3[9]),
    .c(al_eb2b30c3[10]),
    .d(al_eb2b30c3[12]),
    .e(al_eb2b30c3[13]),
    .f(al_eb2b30c3[14]),
    .o(al_35dbcd92));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000100000000))
    al_f6d60342 (
    .a(al_eb2b30c3[1]),
    .b(al_eb2b30c3[2]),
    .c(al_eb2b30c3[4]),
    .d(al_eb2b30c3[5]),
    .e(al_eb2b30c3[6]),
    .f(al_eb2b30c3[7]),
    .o(al_6a936812));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_22c97eef (
    .a(al_35dbcd92),
    .b(al_6a936812),
    .c(al_eb2b30c3[15]),
    .o(al_cc204c06));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_a2f1e76c (
    .a(al_cc204c06),
    .b(al_290af98f),
    .c(al_eb2b30c3[0]),
    .d(al_eb2b30c3[3]),
    .e(al_eb2b30c3[11]),
    .o(al_57b095a8));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_e1a9e385 (
    .a(al_57b095a8),
    .o(al_df9b9d5b[2]));
  AL_DFF_X al_3ea2e640 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e11118e),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_165ae4d7));
  AL_MAP_LUT6 #(
    .EQN("(~(E*~D)*~(F*C*~(B*A)))"),
    .INIT(64'h8f008f8fff00ffff))
    al_6236ba64 (
    .a(al_73bb0740),
    .b(al_496839d3),
    .c(al_26eaf94a),
    .d(al_3f0ffcfa),
    .e(al_e11118e),
    .f(al_d7d3035f),
    .o(al_31ffb8d1));
  AL_MAP_LUT6 #(
    .EQN("~(A*~(E*C*~(~F*~(D*~B))))"),
    .INIT(64'hf5f5555575555555))
    al_950b5fc1 (
    .a(al_31ffb8d1),
    .b(al_7521303d),
    .c(al_faa9857b),
    .d(al_72f63008),
    .e(al_29396e02),
    .f(al_153acd6e),
    .o(al_8e1ef4c5));
  AL_DFF_X al_2400dc0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8e1ef4c5),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_e11118e));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hecb96431))
    al_49e91e0e (
    .a(al_8e143433),
    .b(al_3e1806d9),
    .c(al_5a579dd),
    .d(al_18d64456[0]),
    .e(al_3ac23457[0]),
    .o(al_5743d58d[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_5d503988 (
    .a(al_53f15a3f),
    .b(al_5a579dd),
    .o(al_763891b1));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfdeca8b975642031))
    al_aba57371 (
    .a(al_8e143433),
    .b(al_3e1806d9),
    .c(al_763891b1),
    .d(al_18d64456[0]),
    .e(al_18d64456[1]),
    .f(al_3ac23457[1]),
    .o(al_5743d58d[1]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~((~D*~C))*~(E)+A*~(B)*(~D*~C)*~(E)+~(A)*B*(~D*~C)*~(E)+A*B*(~D*~C)*~(E)+~(A)*~(B)*~((~D*~C))*E+A*~(B)*~((~D*~C))*E+~(A)*B*~((~D*~C))*E+A*B*~((~D*~C))*E+~(A)*~(B)*(~D*~C)*E+~(A)*B*(~D*~C)*E)"),
    .INIT(32'hfff5444e))
    al_6ee570ee (
    .a(al_d0093be6),
    .b(al_618f3df7),
    .c(al_18d64456[0]),
    .d(al_18d64456[1]),
    .e(al_18d64456[2]),
    .o(al_60ceba51));
  AL_MAP_LUT6 #(
    .EQN("(C*~(A*~((~E*D)*~(F)*~(B)+(~E*D)*F*~(B)+~((~E*D))*F*B+(~E*D)*F*B)))"),
    .INIT(64'hd0d0f0d050507050))
    al_997a4563 (
    .a(al_8e143433),
    .b(al_3e1806d9),
    .c(al_60ceba51),
    .d(al_53f15a3f),
    .e(al_5a579dd),
    .f(al_3ac23457[2]),
    .o(al_5743d58d[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_45992ea2 (
    .a(al_d0093be6),
    .b(al_618f3df7),
    .o(al_8e143433));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    al_320f74bf (
    .a(al_d0093be6),
    .b(al_cd3c4af6),
    .c(al_618f3df7),
    .o(al_3e1806d9));
  AL_MAP_LUT6 #(
    .EQN("(E*~A*~(F*~((~D*B))*~(C)+F*(~D*B)*~(C)+~(F)*(~D*B)*C+F*(~D*B)*C))"),
    .INIT(64'h5010000055150000))
    al_9d48d762 (
    .a(al_d0093be6),
    .b(al_53f15a3f),
    .c(al_cd3c4af6),
    .d(al_5a579dd),
    .e(al_618f3df7),
    .f(al_3ac23457[3]),
    .o(al_567c0900));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_c7b24a66 (
    .a(al_18d64456[0]),
    .b(al_18d64456[1]),
    .c(al_18d64456[2]),
    .o(al_ee8c5e52));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~A*~(E@(D*~B))))"),
    .INIT(32'h0e0f0b0a))
    al_77b7f8bf (
    .a(al_8e143433),
    .b(al_3e1806d9),
    .c(al_567c0900),
    .d(al_ee8c5e52),
    .e(al_18d64456[3]),
    .o(al_5743d58d[3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_2a47f6f (
    .a(al_18d64456[0]),
    .b(al_18d64456[1]),
    .c(al_18d64456[2]),
    .d(al_18d64456[3]),
    .o(al_5c754024));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(D)*~(E)*~((F*~C))+A*B*D*~(E)*~((F*~C))+~(A)*~(B)*~(D)*E*~((F*~C))+A*~(B)*~(D)*E*~((F*~C))+~(A)*B*~(D)*E*~((F*~C))+A*~(B)*D*E*~((F*~C))+A*B*~(D)*~(E)*(F*~C)+~(A)*~(B)*D*~(E)*(F*~C)+~(A)*B*D*~(E)*(F*~C)+A*B*D*~(E)*(F*~C)+~(A)*~(B)*~(D)*E*(F*~C)+A*~(B)*~(D)*E*(F*~C)+~(A)*B*~(D)*E*(F*~C)+~(A)*~(B)*D*E*(F*~C)+A*~(B)*D*E*(F*~C)+~(A)*B*D*E*(F*~C))"),
    .INIT(64'h27778d8822778888))
    al_a6157dbf (
    .a(al_d0093be6),
    .b(al_5c754024),
    .c(al_cd3c4af6),
    .d(al_618f3df7),
    .e(al_18d64456[4]),
    .f(al_3ac23457[4]),
    .o(al_5743d58d[4]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~(D)*~(E)*~((F*~C))+A*B*D*~(E)*~((F*~C))+~(A)*~(B)*~(D)*E*~((F*~C))+A*~(B)*~(D)*E*~((F*~C))+~(A)*B*~(D)*E*~((F*~C))+A*~(B)*D*E*~((F*~C))+A*B*~(D)*~(E)*(F*~C)+~(A)*~(B)*D*~(E)*(F*~C)+~(A)*B*D*~(E)*(F*~C)+A*B*D*~(E)*(F*~C)+~(A)*~(B)*~(D)*E*(F*~C)+A*~(B)*~(D)*E*(F*~C)+~(A)*B*~(D)*E*(F*~C)+~(A)*~(B)*D*E*(F*~C)+A*~(B)*D*E*(F*~C)+~(A)*B*D*E*(F*~C))"),
    .INIT(64'h27778d8822778888))
    al_d5c26d4 (
    .a(al_d0093be6),
    .b(al_f5e85a1),
    .c(al_cd3c4af6),
    .d(al_618f3df7),
    .e(al_18d64456[5]),
    .f(al_3ac23457[5]),
    .o(al_5743d58d[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_335acca3 (
    .a(al_cd3c4af6),
    .b(al_3ac23457[6]),
    .o(al_b2d09c6f[6]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*C*D*~((~E*B))*~(F)+A*~(C)*~(D)*(~E*B)*~(F)+A*C*~(D)*(~E*B)*~(F)+A*~(C)*D*(~E*B)*~(F)+~(A)*C*D*(~E*B)*~(F)+A*C*D*(~E*B)*~(F)+~(A)*~(C)*~(D)*~((~E*B))*F+A*~(C)*~(D)*~((~E*B))*F+~(A)*C*~(D)*~((~E*B))*F+A*C*~(D)*~((~E*B))*F+A*~(C)*D*~((~E*B))*F+~(A)*C*D*~((~E*B))*F+A*C*D*~((~E*B))*F+~(A)*~(C)*~(D)*(~E*B)*F+~(A)*C*~(D)*(~E*B)*F+~(A)*C*D*(~E*B)*F)"),
    .INIT(64'hfaff72775000d888))
    al_38533758 (
    .a(al_d0093be6),
    .b(al_f5e85a1),
    .c(al_b2d09c6f[6]),
    .d(al_618f3df7),
    .e(al_18d64456[5]),
    .f(al_18d64456[6]),
    .o(al_5743d58d[6]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_c7dc4a7f (
    .a(al_18d64456[0]),
    .b(al_18d64456[1]),
    .c(al_18d64456[2]),
    .d(al_18d64456[3]),
    .e(al_18d64456[4]),
    .o(al_f5e85a1));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_da0d738d (
    .a(al_f5e85a1),
    .b(al_18d64456[5]),
    .c(al_18d64456[6]),
    .o(al_1520e86d));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*~A))"),
    .INIT(16'h000e))
    al_882fb4 (
    .a(al_72f63008),
    .b(al_153acd6e),
    .c(al_783fafdc),
    .d(al_49948f6),
    .o(al_47214dbf));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~E*~D*~C*A))"),
    .INIT(32'hccccccc4))
    al_82cf35e8 (
    .a(al_f5e85a1),
    .b(al_47214dbf),
    .c(al_18d64456[5]),
    .d(al_18d64456[6]),
    .e(al_18d64456[7]),
    .o(al_d0093be6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(D)*E*~((F*~C))+A*~(B)*~(D)*E*~((F*~C))+~(A)*B*~(D)*E*~((F*~C))+~(A)*B*D*E*~((F*~C))+~(A)*~(B)*D*~(E)*(F*~C)+A*~(B)*D*~(E)*(F*~C)+~(A)*~(B)*~(D)*E*(F*~C)+A*~(B)*~(D)*E*(F*~C)+~(A)*B*~(D)*E*(F*~C)+~(A)*~(B)*D*E*(F*~C)+A*~(B)*D*E*(F*~C)+~(A)*B*D*E*(F*~C))"),
    .INIT(64'h4777030044770000))
    al_20f56ae6 (
    .a(al_1520e86d),
    .b(al_d0093be6),
    .c(al_cd3c4af6),
    .d(al_618f3df7),
    .e(al_18d64456[7]),
    .f(al_3ac23457[7]),
    .o(al_5743d58d[7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_b42865bd (
    .a(al_1520e86d),
    .b(al_153acd6e),
    .c(al_18d64456[7]),
    .o(al_e1b52e50));
  AL_DFF_X al_b2cc10f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1b52e50),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_29396e02));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfef4aaa054540000))
    al_f6802229 (
    .a(al_53f15a3f),
    .b(al_72f63008),
    .c(al_846b6533),
    .d(al_7694b99f),
    .e(al_29396e02),
    .f(al_24faf4d6),
    .o(al_a50584b2));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    al_6852e6d (
    .a(al_b05da9fd),
    .b(al_cd3c4af6),
    .c(al_5a579dd),
    .d(al_7b30ef6a),
    .o(al_c1b27879));
  AL_MAP_LUT6 #(
    .EQN("(~F*~(B*~(C*~(~E*~(~D*A)))))"),
    .INIT(64'h00000000f3f333b3))
    al_74166c2a (
    .a(al_a50584b2),
    .b(al_c1b27879),
    .c(al_7521303d),
    .d(al_6f12ed1d),
    .e(al_153acd6e),
    .f(al_4024362),
    .o(al_160ccdf));
  AL_DFF_X al_f8910726 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_160ccdf),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_b05da9fd));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_12a87508 (
    .a(al_803bd5d9),
    .b(al_1a83737a[0]),
    .c(al_e29488b2[0]),
    .o(al_1d28bc9[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1f5f0e5c (
    .a(al_803bd5d9),
    .b(al_1a83737a[10]),
    .c(al_e29488b2[10]),
    .o(al_1d28bc9[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_24a5fba (
    .a(al_803bd5d9),
    .b(al_1a83737a[11]),
    .c(al_e29488b2[11]),
    .o(al_1d28bc9[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_64b4510a (
    .a(al_803bd5d9),
    .b(al_1a83737a[12]),
    .c(al_e29488b2[12]),
    .o(al_1d28bc9[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c6ba100a (
    .a(al_803bd5d9),
    .b(al_1a83737a[13]),
    .c(al_e29488b2[13]),
    .o(al_1d28bc9[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_eb3b04cb (
    .a(al_803bd5d9),
    .b(al_1a83737a[1]),
    .c(al_e29488b2[1]),
    .o(al_1d28bc9[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8005ea0 (
    .a(al_803bd5d9),
    .b(al_1a83737a[2]),
    .c(al_e29488b2[2]),
    .o(al_1d28bc9[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_575892d9 (
    .a(al_803bd5d9),
    .b(al_1a83737a[3]),
    .c(al_e29488b2[3]),
    .o(al_1d28bc9[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2992bd6f (
    .a(al_803bd5d9),
    .b(al_1a83737a[4]),
    .c(al_e29488b2[4]),
    .o(al_1d28bc9[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ad9c379c (
    .a(al_803bd5d9),
    .b(al_1a83737a[5]),
    .c(al_e29488b2[5]),
    .o(al_1d28bc9[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6f9ad48 (
    .a(al_803bd5d9),
    .b(al_1a83737a[6]),
    .c(al_e29488b2[6]),
    .o(al_1d28bc9[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_de10d141 (
    .a(al_803bd5d9),
    .b(al_1a83737a[7]),
    .c(al_e29488b2[7]),
    .o(al_1d28bc9[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_770e4c88 (
    .a(al_803bd5d9),
    .b(al_1a83737a[8]),
    .c(al_e29488b2[8]),
    .o(al_1d28bc9[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_30ea8167 (
    .a(al_803bd5d9),
    .b(al_1a83737a[9]),
    .c(al_e29488b2[9]),
    .o(al_1d28bc9[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_3ed2863 (
    .a(tx_clk_en),
    .b(al_618f3df7),
    .o(al_86ce862e));
  AL_DFF_X al_fc5c4308 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a231fc3f),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_803bd5d9));
  AL_MAP_LUT5 #(
    .EQN("(~(~C*~B)*~(E*~(~D*A)))"),
    .INIT(32'h00a8fcfc))
    al_8784805c (
    .a(al_7521303d),
    .b(al_72f63008),
    .c(al_846b6533),
    .d(al_b05da9fd),
    .e(al_aaba7825),
    .o(al_f6a2d163));
  AL_MAP_LUT6 #(
    .EQN("(~D*~C*~(~B*~A*~(F*~E)))"),
    .INIT(64'h000e000f000e000e))
    al_b6a67e89 (
    .a(al_f6a2d163),
    .b(al_7694b99f),
    .c(al_7b30ef6a),
    .d(al_153acd6e),
    .e(al_aaba7825),
    .f(al_74608a10),
    .o(al_aa4375dc));
  AL_DFF_X al_d94029f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa4375dc),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3daf6177));
  AL_DFF_X al_79f8fd1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d5178990),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd3c4af6));
  AL_MAP_LUT6 #(
    .EQN("(~B*(E*~(C)*~((~(~F*~D)*A))+E*C*~((~(~F*~D)*A))+~(E)*C*(~(~F*~D)*A)+E*C*(~(~F*~D)*A)))"),
    .INIT(64'h3131202031332000))
    al_7fe17ac7 (
    .a(tx_clk_en),
    .b(al_2dbca608),
    .c(al_5e767b18),
    .d(al_3f0ffcfa),
    .e(al_cd3c4af6),
    .f(al_618f3df7),
    .o(al_d5178990));
  AL_DFF_X al_f25bae5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_46f6a926),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_5ed94f60));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_abd4c9ad (
    .a(al_cae9c79a),
    .b(al_6a6d2547[0]),
    .o(al_2e49f5b3[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_bbe9de6a (
    .a(al_cae9c79a),
    .b(al_6a6d2547[1]),
    .o(al_2e49f5b3[1]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    al_a2068949 (
    .a(al_cae9c79a),
    .b(al_6a6d2547[2]),
    .o(al_2e49f5b3[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_72da748 (
    .a(al_cae9c79a),
    .b(al_6a6d2547[3]),
    .o(al_2e49f5b3[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_16e320c3 (
    .a(al_cae9c79a),
    .b(al_6a6d2547[3]),
    .c(al_6a6d2547[4]),
    .o(al_2e49f5b3[4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(~C*~B)))"),
    .INIT(16'ha802))
    al_f66776b7 (
    .a(al_cae9c79a),
    .b(al_6a6d2547[3]),
    .c(al_6a6d2547[4]),
    .d(al_6a6d2547[5]),
    .o(al_2e49f5b3[5]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(C*~(~B*~A)))"),
    .INIT(32'h0000001f))
    al_850b0c91 (
    .a(al_6a6d2547[0]),
    .b(al_6a6d2547[1]),
    .c(al_6a6d2547[3]),
    .d(al_6a6d2547[6]),
    .e(al_6a6d2547[7]),
    .o(al_66ecf32f));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*~(~E*~D*A))"),
    .INIT(32'h30303010))
    al_1bf2d8b (
    .a(al_66ecf32f),
    .b(al_cd3c4af6),
    .c(al_5ed94f60),
    .d(al_6a6d2547[4]),
    .e(al_6a6d2547[5]),
    .o(al_cae9c79a));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@(~D*~C*~B)))"),
    .INIT(32'haaa80002))
    al_5cc3f1bb (
    .a(al_cae9c79a),
    .b(al_6a6d2547[3]),
    .c(al_6a6d2547[4]),
    .d(al_6a6d2547[5]),
    .e(al_6a6d2547[6]),
    .o(al_2e49f5b3[6]));
  AL_MAP_LUT6 #(
    .EQN("(F*A*~(~E*~D*~C*~B))"),
    .INIT(64'haaaaaaa800000000))
    al_27689259 (
    .a(al_cae9c79a),
    .b(al_6a6d2547[3]),
    .c(al_6a6d2547[4]),
    .d(al_6a6d2547[5]),
    .e(al_6a6d2547[6]),
    .f(al_6a6d2547[7]),
    .o(al_2e49f5b3[7]));
  AL_DFF_X al_d121ad10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1ea4ba5b),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_db1fbb11));
  AL_DFF_X al_e511d66a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6b8a9b19),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_55ac2d11));
  AL_DFF_X al_cb7eeacf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_75707d25),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d1cfb12d));
  AL_DFF_X al_133f6b2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_de9cd38),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_5a579dd));
  AL_DFF_X al_9db00c23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f396fdd4),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_5c82d563));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    al_4053b3f3 (
    .a(al_cc204c06),
    .b(al_eb2b30c3[0]),
    .c(al_eb2b30c3[3]),
    .d(al_eb2b30c3[11]),
    .o(al_a2faab7b));
  AL_DFF_X al_e3b11705 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9a990f97),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f12ed1d));
  AL_MAP_LUT6 #(
    .EQN("(~C*(D*~((~E*A))*~((F*B))+D*(~E*A)*~((F*B))+~(D)*(~E*A)*(F*B)+D*(~E*A)*(F*B)))"),
    .INIT(64'h03000b080f000f00))
    al_c02977aa (
    .a(al_73bb0740),
    .b(tx_clk_en),
    .c(al_2dbca608),
    .d(al_6f12ed1d),
    .e(al_2162c82e),
    .f(al_4024362),
    .o(al_9a990f97));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~C)*~(D*~B*A))"),
    .INIT(32'hddffd0f0))
    al_8b3e3520 (
    .a(al_ff9a0466),
    .b(al_53f15a3f),
    .c(al_9b760ae7),
    .d(al_618f3df7),
    .e(al_34e054a0),
    .o(al_14c1cb65));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    al_29cc7876 (
    .a(al_b241735d),
    .b(al_14c1cb65),
    .c(al_bfd01551),
    .o(al_290f1a7e));
  AL_DFF_X al_2156eaa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_290f1a7e),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_9b760ae7));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h88a0))
    al_b6ffa4f0 (
    .a(al_cd3c4af6),
    .b(al_9b760ae7),
    .c(al_ef80f5cf),
    .d(al_4024362),
    .o(al_32e957a5));
  AL_DFF_X al_6919e46a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_32e957a5),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_ef80f5cf));
  AL_MAP_LUT5 #(
    .EQN("~(~(~D*B)*~(~E*C*A))"),
    .INIT(32'h00cca0ec))
    al_fe8fc269 (
    .a(al_cf20ff1a),
    .b(al_d8c8c74d),
    .c(al_7b30ef6a),
    .d(al_34e054a0),
    .e(al_c9168fb8[5]),
    .o(al_36c5508));
  AL_DFF_X al_2c379876 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_36c5508),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d8c8c74d));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*B)*~(~C*A))"),
    .INIT(16'h0ace))
    al_65417374 (
    .a(al_5dda436f),
    .b(al_96ecb37f),
    .c(al_34e054a0),
    .d(al_b4f442b4),
    .o(al_c6a375ec));
  AL_DFF_X al_777c841a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c6a375ec),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_5dda436f));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_11a8e72a (
    .a(al_4bdde34),
    .b(al_136addab),
    .c(al_c9c0fa32),
    .d(al_8e6107a7),
    .e(al_15bf91ee),
    .f(al_af4842d7),
    .o(al_3e1dba29));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_33178e63 (
    .a(al_3e1dba29),
    .b(al_336bd542),
    .o(al_71ed2e0a));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~B)*~(~C*A))"),
    .INIT(16'h3b0a))
    al_99f13b36 (
    .a(al_78612548),
    .b(al_2c24255b),
    .c(al_618f3df7),
    .d(al_b4f442b4),
    .o(al_64320b18));
  AL_DFF_X al_bd01fd8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64320b18),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_78612548));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(A*~(~E*~D*~B)))"),
    .INIT(32'h05050507))
    al_c63d85bb (
    .a(al_adc2de29),
    .b(al_c8a3ac58),
    .c(al_2c24255b),
    .d(al_618f3df7),
    .e(al_4024362),
    .o(al_46d73024));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_cc4a2224 (
    .a(al_46d73024),
    .b(al_5c82d563),
    .c(al_34e054a0),
    .o(al_4ce1f25a));
  AL_DFF_X al_9840d6eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4ce1f25a),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2c24255b));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(~C*~A))"),
    .INIT(16'h0032))
    al_d7b740f7 (
    .a(al_adc2de29),
    .b(al_5c82d563),
    .c(al_2162c82e),
    .d(al_34e054a0),
    .o(al_b02bbd88));
  AL_DFF_X al_5b930d31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b02bbd88),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2162c82e));
  AL_DFF_X al_b2a730c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b1d9ebd5),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_290af98f));
  AL_MAP_LUT3 #(
    .EQN("~(A*(C@B))"),
    .INIT(8'hd7))
    al_274e1540 (
    .a(al_7b30ef6a),
    .b(al_3ab98f26[0]),
    .c(al_3ab98f26[1]),
    .o(al_9bde74c4[1]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(~E*~(C*~(B*~A))))"),
    .INIT(32'hff00b000))
    al_151eed6a (
    .a(al_3fc75a33),
    .b(al_a8e6ffb8),
    .c(al_35f24fff),
    .d(al_ac79ddb),
    .e(al_7b30ef6a),
    .o(al_870286f7));
  AL_DFF_X al_476c2a1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_870286f7),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_7b30ef6a));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_4a16657d (
    .a(al_e101ff9a),
    .b(al_7dd23876),
    .o(al_adc2de29));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_e94be992 (
    .a(al_b241735d),
    .b(al_72f63008),
    .c(al_e9ae3746),
    .o(al_a8e6ffb8));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_e60e26cb (
    .a(al_efdbdafe),
    .b(al_e11118e),
    .o(al_35f24fff));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_7283de3e (
    .a(al_3f0ffcfa),
    .b(al_153acd6e),
    .c(al_49948f6),
    .d(al_d7d3035f),
    .o(al_ac79ddb));
  AL_MAP_LUT6 #(
    .EQN("(D*(E*~(F)*~((C*~(B*~A)))+E*F*~((C*~(B*~A)))+~(E)*F*(C*~(B*~A))+E*F*(C*~(B*~A))))"),
    .INIT(64'hff00b0004f000000))
    al_1314006d (
    .a(al_3fc75a33),
    .b(al_a8e6ffb8),
    .c(al_35f24fff),
    .d(al_ac79ddb),
    .e(al_96ecb37f),
    .f(al_ebd2d7),
    .o(al_482b5978));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_c3c81ba7 (
    .a(al_2a1554ab[0]),
    .b(al_2a1554ab[1]),
    .c(al_2a1554ab[2]),
    .o(al_da48a386));
  AL_MAP_LUT6 #(
    .EQN("(~C*~(~E*~D*~(~A*~(~F*~B))))"),
    .INIT(64'h0f0f0f050f0f0f04))
    al_c785fe44 (
    .a(al_b5c79ef6),
    .b(al_9ba351db),
    .c(al_7b30ef6a),
    .d(al_2d5ca5c8),
    .e(al_cb8cffb4[2]),
    .f(al_931288d8[1]),
    .o(al_b241735d));
  AL_MAP_LUT6 #(
    .EQN("(~(~(E*C)*~(~D*B))*~(~F*~A))"),
    .INIT(64'hf0fc00cca0a80088))
    al_db7700c0 (
    .a(al_da48a386),
    .b(al_adc2de29),
    .c(al_266f6c4c),
    .d(al_7b30ef6a),
    .e(al_6b8a9b19),
    .f(al_4024362),
    .o(al_e5994b5e));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~E*D*~C*~A))"),
    .INIT(32'h33333233))
    al_733c20ec (
    .a(al_53f15a3f),
    .b(al_3daf6177),
    .c(al_d1cfb12d),
    .d(al_9953d0c8),
    .e(al_cb8cffb4[2]),
    .o(al_a2667927));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_a15e22a1 (
    .a(al_e5994b5e),
    .b(al_a2667927),
    .o(al_3fc75a33));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(~C*~B))"),
    .INIT(16'h00a8))
    al_b9cba1ce (
    .a(al_cd3c4af6),
    .b(al_fb660f65),
    .c(al_f65615d7),
    .d(al_cb8cffb4[1]),
    .o(al_efdbdafe));
  AL_DFF_X al_4b3129b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_482b5978),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_96ecb37f));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_e4280332 (
    .a(al_9e425de4),
    .b(al_3ce55a07[0]),
    .o(al_2e44f12e[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    al_ba0e9785 (
    .a(al_9e425de4),
    .b(al_3ce55a07[0]),
    .c(al_3ce55a07[1]),
    .o(al_2e44f12e[1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(C*B)))"),
    .INIT(16'h2a80))
    al_55f9b050 (
    .a(al_9e425de4),
    .b(al_3ce55a07[0]),
    .c(al_3ce55a07[1]),
    .d(al_3ce55a07[2]),
    .o(al_2e44f12e[2]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@(D*C*B)))"),
    .INIT(32'h2aaa8000))
    al_5a318338 (
    .a(al_9e425de4),
    .b(al_3ce55a07[0]),
    .c(al_3ce55a07[1]),
    .d(al_3ce55a07[2]),
    .e(al_3ce55a07[3]),
    .o(al_2e44f12e[3]));
  AL_MAP_LUT6 #(
    .EQN("(A*(F@(E*D*C*B)))"),
    .INIT(64'h2aaaaaaa80000000))
    al_286714f8 (
    .a(al_9e425de4),
    .b(al_3ce55a07[0]),
    .c(al_3ce55a07[1]),
    .d(al_3ce55a07[2]),
    .e(al_3ce55a07[3]),
    .f(al_3ce55a07[4]),
    .o(al_2e44f12e[4]));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_91b93e2e (
    .a(al_3ce55a07[0]),
    .b(al_3ce55a07[1]),
    .c(al_3ce55a07[2]),
    .d(al_3ce55a07[3]),
    .e(al_3ce55a07[4]),
    .f(al_3ce55a07[5]),
    .o(al_302a167b[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_4859d44e (
    .a(al_9e425de4),
    .b(al_302a167b[5]),
    .o(al_2e44f12e[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    al_1eb65662 (
    .a(al_9e425de4),
    .b(al_a7784e58),
    .c(al_3ce55a07[6]),
    .o(al_2e44f12e[6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(C*B)))"),
    .INIT(16'h2a80))
    al_68895f86 (
    .a(al_9e425de4),
    .b(al_a7784e58),
    .c(al_3ce55a07[6]),
    .d(al_3ce55a07[7]),
    .o(al_2e44f12e[7]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@(D*C*B)))"),
    .INIT(32'h2aaa8000))
    al_e040c35f (
    .a(al_9e425de4),
    .b(al_a7784e58),
    .c(al_3ce55a07[6]),
    .d(al_3ce55a07[7]),
    .e(al_3ce55a07[8]),
    .o(al_2e44f12e[8]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_f93afdc5 (
    .a(al_3ce55a07[0]),
    .b(al_3ce55a07[1]),
    .c(al_3ce55a07[2]),
    .d(al_3ce55a07[3]),
    .e(al_3ce55a07[4]),
    .f(al_3ce55a07[5]),
    .o(al_a7784e58));
  AL_MAP_LUT6 #(
    .EQN("(A*(F@(E*D*C*B)))"),
    .INIT(64'h2aaaaaaa80000000))
    al_f86a2506 (
    .a(al_9e425de4),
    .b(al_a7784e58),
    .c(al_3ce55a07[6]),
    .d(al_3ce55a07[7]),
    .e(al_3ce55a07[8]),
    .f(al_3ce55a07[9]),
    .o(al_2e44f12e[9]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_c57afc8 (
    .a(al_ff9a0466),
    .b(al_cd3c4af6),
    .c(al_5a579dd),
    .o(al_7521303d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_551fb681 (
    .a(al_3ce55a07[0]),
    .b(al_3ce55a07[1]),
    .c(al_3ce55a07[2]),
    .d(al_3ce55a07[3]),
    .e(al_3ce55a07[4]),
    .f(al_3ce55a07[5]),
    .o(al_37168961));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_1550e3ab (
    .a(al_37168961),
    .b(al_efdbdafe),
    .c(al_3ce55a07[7]),
    .d(al_3ce55a07[8]),
    .o(al_b48e2d4e));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(A*(B*D*~(E)+~(B)*~(D)*E)))"),
    .INIT(32'h0f0d070f))
    al_7f1e11ff (
    .a(al_b48e2d4e),
    .b(al_5a579dd),
    .c(al_ebd2d7),
    .d(al_3ce55a07[6]),
    .e(al_3ce55a07[9]),
    .o(al_efc518d8));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(~C*B)))"),
    .INIT(16'h0455))
    al_c7a4f022 (
    .a(al_efc518d8),
    .b(al_7521303d),
    .c(al_53f15a3f),
    .d(al_618f3df7),
    .o(al_857e17ab));
  AL_DFF_X al_d1aff26f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_857e17ab),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_ebd2d7));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*C*~B*A)"),
    .INIT(64'h0000000000000020))
    al_4fcb3bb7 (
    .a(al_5305cb61[8]),
    .b(al_5305cb61[9]),
    .c(al_5305cb61[10]),
    .d(al_5305cb61[11]),
    .e(al_5305cb61[12]),
    .f(al_5305cb61[13]),
    .o(al_5ce38362));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*~B*~A)"),
    .INIT(64'h1000000000000000))
    al_3671fbb0 (
    .a(al_153acd6e),
    .b(al_5305cb61[0]),
    .c(al_5305cb61[1]),
    .d(al_5305cb61[5]),
    .e(al_5305cb61[6]),
    .f(al_5305cb61[7]),
    .o(al_e0dc1ae0));
  AL_MAP_LUT4 #(
    .EQN("(~C*(~(A)*~(B)*~(D)+A*B*D))"),
    .INIT(16'h0801))
    al_41cf5310 (
    .a(al_5305cb61[2]),
    .b(al_5305cb61[3]),
    .c(al_5305cb61[14]),
    .d(al_e31e36f5[2]),
    .o(al_762c3367));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    al_de2cb788 (
    .a(al_5ce38362),
    .b(al_e0dc1ae0),
    .c(al_762c3367),
    .d(al_58e1cc88),
    .e(al_5305cb61[4]),
    .o(al_dcbb090f));
  AL_MAP_LUT6 #(
    .EQN("(~D*~(~A*~(E*~(C*~(~F*~B)))))"),
    .INIT(64'h00af00aa00bf00aa))
    al_bcb92a59 (
    .a(al_dcbb090f),
    .b(al_72f63008),
    .c(al_29396e02),
    .d(al_db1fbb11),
    .e(al_6b8a9b19),
    .f(al_153acd6e),
    .o(al_67b72f88));
  AL_DFF_X al_8dfe5e67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_67b72f88),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_6b8a9b19));
  AL_MAP_LUT6 #(
    .EQN("(B*~(~(~F*C)*~(D*~(E*~A))))"),
    .INIT(64'h8800cc00c8c0ccc0))
    al_157f4e7f (
    .a(al_efdbdafe),
    .b(al_7521303d),
    .c(al_53f15a3f),
    .d(al_6f12ed1d),
    .e(al_2162c82e),
    .f(al_24faf4d6),
    .o(al_aa32962e));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(C*~B)*~(E*~A))"),
    .INIT(32'hff75ff30))
    al_726eee0d (
    .a(al_aa32962e),
    .b(al_e11118e),
    .c(al_153acd6e),
    .d(al_49948f6),
    .e(al_b4f442b4),
    .o(al_94871a17));
  AL_DFF_X al_95946742 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_94871a17),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_153acd6e));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(~B*A))"),
    .INIT(8'hf2))
    al_8129c801 (
    .a(al_b96742e9),
    .b(al_618f3df7),
    .c(al_5305cb61[6]),
    .o(al_6f78b0c1));
  AL_DFF_X al_cd9185dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6f78b0c1),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_b96742e9));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*~A)"),
    .INIT(32'h00000010))
    al_be0c6265 (
    .a(al_3f0ffcfa),
    .b(al_e11118e),
    .c(al_cd3c4af6),
    .d(al_5a579dd),
    .e(al_7b30ef6a),
    .o(al_8a331b5c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_a8894927 (
    .a(al_1b8c3389[3]),
    .b(al_1b8c3389[4]),
    .c(al_1b8c3389[5]),
    .d(al_1b8c3389[6]),
    .e(al_1b8c3389[7]),
    .f(al_1b8c3389[8]),
    .o(al_76e16a6c));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~(A*~(C*B))))"),
    .INIT(32'h00002aff))
    al_23fb1ad1 (
    .a(al_76e16a6c),
    .b(al_1b8c3389[1]),
    .c(al_1b8c3389[2]),
    .d(al_1b8c3389[9]),
    .e(al_1b8c3389[10]),
    .o(al_3fe47357));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~A*~(D*~C*~B)))"),
    .INIT(32'h0000abaa))
    al_77eea98b (
    .a(al_3fe47357),
    .b(al_e5994b5e),
    .c(al_b241735d),
    .d(al_a2667927),
    .e(al_aaba7825),
    .o(al_250851df));
  AL_MAP_LUT4 #(
    .EQN("~(~D*C*~(B*~A))"),
    .INIT(16'hff4f))
    al_ad400d45 (
    .a(al_250851df),
    .b(al_8a331b5c),
    .c(al_cd3c4af6),
    .d(al_5a579dd),
    .o(al_63eeda3d));
  AL_DFF_X al_53d298b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_63eeda3d),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_aaba7825));
  AL_DFF_X al_b11936f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f5fd4d02),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2d5ca5c8));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_31983773 (
    .a(al_f8ee3a1f),
    .b(al_8c6e2d36),
    .o(al_765cb78c));
  AL_DFF_X al_ffb05bb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_765cb78c),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f5fd4d02));
  AL_DFF_X al_56a43ede (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3bac4202),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_9953d0c8));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    al_517dbe7d (
    .a(al_618f3df7),
    .b(al_2a1554ab[0]),
    .o(al_cf2a0a44[0]));
  AL_MAP_LUT3 #(
    .EQN("~(A*(C@B))"),
    .INIT(8'hd7))
    al_6d7bff3e (
    .a(al_618f3df7),
    .b(al_2a1554ab[0]),
    .c(al_2a1554ab[1]),
    .o(al_cf2a0a44[1]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(D@(~C*~B)))"),
    .INIT(16'hfd57))
    al_85c7f80d (
    .a(al_618f3df7),
    .b(al_2a1554ab[0]),
    .c(al_2a1554ab[1]),
    .d(al_2a1554ab[2]),
    .o(al_cf2a0a44[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_1a68c8ed (
    .a(al_618f3df7),
    .b(al_4024362),
    .o(al_3bac4202));
  AL_MAP_LUT5 #(
    .EQN("(D*~(~E*~C*~(~B*~A)))"),
    .INIT(32'hff00f100))
    al_9bb18139 (
    .a(al_fff0fd72[0]),
    .b(al_fff0fd72[1]),
    .c(al_fff0fd72[2]),
    .d(al_3f0ffcfa),
    .e(al_130ad14e),
    .o(al_8c59fe48));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(~F*~(~C*~(E*D*B))))"),
    .INIT(64'haaaaaaaafefafafa))
    al_cb015858 (
    .a(al_8c59fe48),
    .b(al_7521303d),
    .c(al_3bac4202),
    .d(al_72f63008),
    .e(al_29396e02),
    .f(al_7b30ef6a),
    .o(al_27722f64));
  AL_DFF_X al_ccc238a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_27722f64),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618f3df7));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    al_16ab761c (
    .a(al_9953d0c8),
    .b(al_2a1554ab[0]),
    .c(al_2a1554ab[1]),
    .d(al_2a1554ab[2]),
    .o(al_388a24e));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*C*~(D)*~((~E*B))+A*C*~(D)*~((~E*B))+~(A)*C*D*~((~E*B))+~(A)*~(C)*~(D)*(~E*B)+A*~(C)*~(D)*(~E*B)+~(A)*C*~(D)*(~E*B)+A*C*~(D)*(~E*B))"),
    .INIT(32'h50f010fc))
    al_e778a6 (
    .a(al_388a24e),
    .b(al_73bb0740),
    .c(al_bfd01551),
    .d(al_c0e7d6fc),
    .e(al_a381b363),
    .o(al_fb3b1f47));
  AL_DFF_X al_98cda960 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_fb3b1f47),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_bfd01551));
  AL_DFF_X al_29052d5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(gmii_col),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_fb660f65));
  AL_DFF_X al_3aedad3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4e287126),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_c0e7d6fc));
  AL_DFF_X al_242ec5bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_73bb0740),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_a381b363));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_20bcea04 (
    .a(al_59a6ee8e[8]),
    .b(al_59a6ee8e[9]),
    .c(al_59a6ee8e[10]),
    .d(al_59a6ee8e[11]),
    .e(al_59a6ee8e[12]),
    .f(al_59a6ee8e[13]),
    .o(al_de2d167c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_d777e001 (
    .a(al_59a6ee8e[2]),
    .b(al_59a6ee8e[3]),
    .c(al_59a6ee8e[4]),
    .d(al_59a6ee8e[5]),
    .e(al_59a6ee8e[6]),
    .f(al_59a6ee8e[7]),
    .o(al_da5e606a));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_2d552337 (
    .a(al_de2d167c),
    .b(al_da5e606a),
    .c(al_59a6ee8e[0]),
    .d(al_59a6ee8e[1]),
    .e(al_59a6ee8e[14]),
    .o(al_f5fb13b0));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(~C*B))"),
    .INIT(8'hae))
    al_d3487a9e (
    .a(al_f5fb13b0),
    .b(al_84db8eae),
    .c(al_34e054a0),
    .o(al_27b5418b));
  AL_DFF_X al_fe50d69e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_27b5418b),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_84db8eae));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~F*~E)*~((~B*~A))*~(D)+(~F*~E)*(~B*~A)*~(D)+~((~F*~E))*(~B*~A)*D+(~F*~E)*(~B*~A)*D))"),
    .INIT(64'he0f0e0f0e0f0e000))
    al_8a1a394e (
    .a(al_d32c67d0),
    .b(al_31529785),
    .c(al_cd3c4af6),
    .d(al_5a579dd),
    .e(al_62aa372c),
    .f(al_6ed289d3),
    .o(al_9e425de4));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    al_452b538d (
    .a(al_cd3c4af6),
    .b(al_7b30ef6a),
    .c(al_f65615d7),
    .d(al_d7d3035f),
    .o(al_f3e72725));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*B)*~(D*~(~C*~A)))"),
    .INIT(32'hfeccfa00))
    al_6d86846b (
    .a(al_3fc75a33),
    .b(al_9e425de4),
    .c(al_b241735d),
    .d(al_f3e72725),
    .e(al_fb660f65),
    .o(al_fe5b64db));
  AL_DFF_X al_e53051a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_fe5b64db),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f65615d7));
  AL_DFF_X al_34d4b2df (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_da48a386),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1717406d));
  AL_DFF_X al_1502ae0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9953d0c8),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cd9f7a57));
  AL_DFF_X al_907cb524 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e9ae3746),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_74608a10));
  AL_MAP_LUT5 #(
    .EQN("(~E*C*A*~(~D*~B))"),
    .INIT(32'h0000a080))
    al_51b7cf9b (
    .a(al_faa9857b),
    .b(al_72f63008),
    .c(al_29396e02),
    .d(al_153acd6e),
    .e(al_34e054a0),
    .o(al_a78f40cd));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(~E*D*~C*B))"),
    .INIT(32'haaaaaeaa))
    al_4816c261 (
    .a(al_a78f40cd),
    .b(al_cd3c4af6),
    .c(al_5a579dd),
    .d(al_34e054a0),
    .e(al_4024362),
    .o(al_a3d91059));
  AL_DFF_X al_19c8dbb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3d91059),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_34e054a0));
  AL_DFF_X al_2b4c8c36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a2faab7b),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_862844a1));
  AL_DFF_X al_82f722bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d32c67d0),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_62aa372c));
  AL_DFF_X al_67858766 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_31529785),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_6ed289d3));
  AL_DFF_X al_6e67242a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_57b095a8),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_58e1cc88));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*~A)"),
    .INIT(32'h00000010))
    al_65a6cb14 (
    .a(al_e11118e),
    .b(al_7b30ef6a),
    .c(al_e9ae3746),
    .d(al_49948f6),
    .e(al_b4f442b4),
    .o(al_7c0f8e52));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(~(~D*~(F*C))*~(B)*~(E)+~(~D*~(F*C))*B*~(E)+~(~(~D*~(F*C)))*B*E+~(~D*~(F*C))*B*E))"),
    .INIT(64'heeeefffaeeeeffaa))
    al_e4a71cfd (
    .a(al_7c0f8e52),
    .b(al_376757cc),
    .c(al_8c6e2d36),
    .d(al_266f6c4c),
    .e(al_803bd5d9),
    .f(al_b96742e9),
    .o(al_4a2b9f40));
  AL_DFF_X al_54c330e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4a2b9f40),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e9ae3746));
  AL_MAP_LUT5 #(
    .EQN("~(~(C*~B)*~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))"),
    .INIT(32'hff75ba30))
    al_6b1ec69f (
    .a(al_5a579dd),
    .b(al_618f3df7),
    .c(al_24faf4d6),
    .d(al_5305cb61[6]),
    .e(al_5305cb61[9]),
    .o(al_5c9e751b));
  AL_DFF_X al_c0111ecc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5c9e751b),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_24faf4d6));
  AL_DFF_X al_8e2949de (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a78f40cd),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vld));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    al_57ef5311 (
    .a(al_6b8a9b19),
    .b(al_618f3df7),
    .c(al_26e8cb8e),
    .o(al_abe786cc));
  AL_DFF_X al_cd2a889d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_abe786cc),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_26e8cb8e));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    al_92b8a07d (
    .a(al_8c6e2d36),
    .b(al_266f6c4c),
    .c(al_9ba351db),
    .d(al_618f3df7),
    .e(al_4024362),
    .o(al_b1649623));
  AL_DFF_X al_8bae0dea (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b1649623),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_bd8e6c56));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_1d86a3b7 (
    .a(al_7f4e8532),
    .b(al_12ae2ff1),
    .c(al_49948f6),
    .o(al_a3ff8a2f));
  AL_DFF_X al_4ce6c10f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a3ff8a2f),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_783fafdc));
  AL_DFF_X al_372d0e12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49948f6),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_7f4e8532));
  AL_DFF_X al_6a32b8c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7f4e8532),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_12ae2ff1));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_be67fce (
    .a(al_7b30ef6a),
    .b(al_3ab98f26[0]),
    .o(al_9bde74c4[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_a22d8867 (
    .a(al_9bde74c4[0]),
    .b(al_3ab98f26[1]),
    .o(al_f396fdd4));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~C*~(~D*B)))"),
    .INIT(16'ha0a8))
    al_b2079eb4 (
    .a(al_f396fdd4),
    .b(al_cf20ff1a),
    .c(al_96ecb37f),
    .d(al_c9168fb8[5]),
    .o(al_bdf8d79f));
  AL_MAP_LUT6 #(
    .EQN("(D*((F*~(C*B))*~(A)*~(E)+(F*~(C*B))*A*~(E)+~((F*~(C*B)))*A*E+(F*~(C*B))*A*E))"),
    .INIT(64'haa003f00aa000000))
    al_21bb63f4 (
    .a(al_31529785),
    .b(al_ff9a0466),
    .c(al_9aa134ca),
    .d(al_cd3c4af6),
    .e(al_5a579dd),
    .f(al_6ed289d3),
    .o(al_f07e3782));
  AL_MAP_LUT6 #(
    .EQN("(~C*B*~(D*(F*~(A)*~(E)+F*A*~(E)+~(F)*A*E+F*A*E)))"),
    .INIT(64'h040c000c040c0c0c))
    al_f1c81e37 (
    .a(al_d32c67d0),
    .b(al_f718b05a),
    .c(al_3d294c28),
    .d(al_cd3c4af6),
    .e(al_5a579dd),
    .f(al_62aa372c),
    .o(al_6d77788f));
  AL_MAP_LUT6 #(
    .EQN("(~D*~(~F*~A*~(E*C*~B)))"),
    .INIT(64'h00ff00ff00ba00aa))
    al_e693594d (
    .a(al_bdf8d79f),
    .b(al_f07e3782),
    .c(al_6d77788f),
    .d(al_153acd6e),
    .e(al_e9ae3746),
    .f(al_49948f6),
    .o(al_f2f998df));
  AL_DFF_X al_b15a2e45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f2f998df),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_49948f6));
  AL_MAP_LUT6 #(
    .EQN("(F*~D*~(B*(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)))"),
    .INIT(64'h0073007f00000000))
    al_fca63dd6 (
    .a(al_d32c67d0),
    .b(al_cd3c4af6),
    .c(al_5a579dd),
    .d(al_7b30ef6a),
    .e(al_62aa372c),
    .f(al_e9ae3746),
    .o(al_232d54d1));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    al_645b753e (
    .a(al_72f63008),
    .b(al_7694b99f),
    .c(al_7b30ef6a),
    .d(al_153acd6e),
    .e(al_b4f442b4),
    .o(al_465185e7));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(E*~D*~C*A))"),
    .INIT(32'hcccecccc))
    al_2d158175 (
    .a(al_232d54d1),
    .b(al_465185e7),
    .c(al_efdbdafe),
    .d(al_f718b05a),
    .e(al_3d294c28),
    .o(al_4c288bd1));
  AL_DFF_X al_cc5f416c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4c288bd1),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_b4f442b4));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    al_87a6e745 (
    .a(al_3f0ffcfa),
    .b(al_8c6e2d36),
    .c(al_266f6c4c),
    .d(al_7b30ef6a),
    .e(al_4024362),
    .o(al_ec82248c));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    al_3f0068cb (
    .a(al_ec82248c),
    .b(al_da48a386),
    .c(al_618f3df7),
    .o(al_11d61e7f));
  AL_DFF_X al_53bb5b88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_11d61e7f),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_4024362));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~E*D*~B*~A))"),
    .INIT(32'h0f0f0e0f))
    al_2411cdf6 (
    .a(al_165ae4d7),
    .b(al_7b30ef6a),
    .c(al_618f3df7),
    .d(al_130ad14e),
    .e(al_d7d3035f),
    .o(al_32e05e5d));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_b9bddf9c (
    .a(al_32e05e5d),
    .b(al_cd3c4af6),
    .c(al_5a579dd),
    .o(al_e9c121e6));
  AL_DFF_X al_402bd109 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e9c121e6),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_130ad14e));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(~D*B))"),
    .INIT(16'h0a02))
    al_47f9f59c (
    .a(al_f396fdd4),
    .b(al_cf20ff1a),
    .c(al_96ecb37f),
    .d(al_c9168fb8[5]),
    .o(al_75707d25));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~D*~C*~B))"),
    .INIT(32'haaabaaaa))
    al_48b3a5ea (
    .a(al_75707d25),
    .b(al_3f0ffcfa),
    .c(al_e11118e),
    .d(al_153acd6e),
    .e(al_d7d3035f),
    .o(al_571ce91a));
  AL_DFF_X al_e51a0192 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_571ce91a),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d7d3035f));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_b8e313d5 (
    .a(1'b0),
    .o({al_968a4ecb,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6fb5d77f (
    .a(al_5305cb61[0]),
    .b(1'b1),
    .c(al_968a4ecb),
    .o({al_26e81f34,al_b7d1cff2[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b8a1df91 (
    .a(al_5305cb61[1]),
    .b(1'b0),
    .c(al_26e81f34),
    .o({al_9ea76e6c,al_b7d1cff2[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b6c03793 (
    .a(al_5305cb61[2]),
    .b(1'b0),
    .c(al_9ea76e6c),
    .o({al_63060b04,al_b7d1cff2[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9304f7c7 (
    .a(al_5305cb61[3]),
    .b(1'b0),
    .c(al_63060b04),
    .o({al_3171227d,al_b7d1cff2[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d7e21145 (
    .a(al_5305cb61[4]),
    .b(1'b0),
    .c(al_3171227d),
    .o({al_360de72,al_b7d1cff2[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c3d4fffb (
    .a(al_5305cb61[5]),
    .b(1'b0),
    .c(al_360de72),
    .o({al_e707cc0b,al_b7d1cff2[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_609fe06b (
    .a(al_5305cb61[6]),
    .b(1'b0),
    .c(al_e707cc0b),
    .o({al_84db4232,al_b7d1cff2[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b3d6899f (
    .a(al_5305cb61[7]),
    .b(1'b0),
    .c(al_84db4232),
    .o({al_6a7aee90,al_b7d1cff2[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_155c05aa (
    .a(al_5305cb61[8]),
    .b(1'b0),
    .c(al_6a7aee90),
    .o({al_af35a257,al_b7d1cff2[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_50c59fe6 (
    .a(al_5305cb61[9]),
    .b(1'b0),
    .c(al_af35a257),
    .o({al_7fda34f5,al_b7d1cff2[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fe5dbeda (
    .a(al_5305cb61[10]),
    .b(1'b0),
    .c(al_7fda34f5),
    .o({al_318f23df,al_b7d1cff2[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3c70ee92 (
    .a(al_5305cb61[11]),
    .b(1'b0),
    .c(al_318f23df),
    .o({al_8202a39,al_b7d1cff2[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_32f0fdfe (
    .a(al_5305cb61[12]),
    .b(1'b0),
    .c(al_8202a39),
    .o({al_33069608,al_b7d1cff2[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ddaa6af1 (
    .a(al_5305cb61[13]),
    .b(1'b0),
    .c(al_33069608),
    .o({al_b430139c,al_b7d1cff2[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1fab4ad9 (
    .a(al_5305cb61[14]),
    .b(1'b0),
    .c(al_b430139c),
    .o({open_n15,al_b7d1cff2[14]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_618f1c1b (
    .a(tx_clk_en),
    .b(al_72f63008),
    .c(al_7694b99f),
    .d(al_c8a3ac58),
    .e(al_7b30ef6a),
    .f(al_153acd6e),
    .o(al_e7b257ab));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_edee51a9 (
    .a(al_e7b257ab),
    .b(al_74608a10),
    .o(al_5ce3a1c4));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_3a98f72a (
    .a(tx_clk_en),
    .b(al_cb8cffb4[13]),
    .o(al_221dcc8d));
  AL_DFF_X al_7886323c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_55a9d56d[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_c9168fb8[0]));
  AL_DFF_X al_678201e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_55a9d56d[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_c9168fb8[1]));
  AL_DFF_X al_f684356f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_55a9d56d[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_c9168fb8[2]));
  AL_DFF_X al_ee7b651e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_55a9d56d[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_c9168fb8[3]));
  AL_DFF_X al_ee3de878 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_55a9d56d[4]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_c9168fb8[4]));
  AL_DFF_X al_37b78ee7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_55a9d56d[5]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_c9168fb8[5]));
  AL_DFF_X al_c5972fae (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[8]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[8]));
  AL_DFF_X al_841a19ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[9]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[9]));
  AL_DFF_X al_d7f93560 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[10]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[10]));
  AL_DFF_X al_4e0d8c38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[0]));
  AL_DFF_X al_106fadcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[1]));
  AL_DFF_X al_dd186eae (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[2]));
  AL_DFF_X al_14ce66ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[3]));
  AL_DFF_X al_46f70bde (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[4]));
  AL_DFF_X al_d010c8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[5]));
  AL_DFF_X al_f0430569 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[6]));
  AL_DFF_X al_d52e1daa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee979a13[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1b8c3389[7]));
  AL_DFF_X al_9caf5efb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[8]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[8]));
  AL_DFF_X al_6cfd8d91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[9]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[9]));
  AL_DFF_X al_2de09edd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[10]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[10]));
  AL_DFF_X al_63532c82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[11]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[11]));
  AL_DFF_X al_ae5adb6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[12]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[12]));
  AL_DFF_X al_a876d3de (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[13]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[13]));
  AL_DFF_X al_98e5956c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[14]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[14]));
  AL_DFF_X al_e2a8a99f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[0]));
  AL_DFF_X al_2320aad5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[1]));
  AL_DFF_X al_6e399b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[2]));
  AL_DFF_X al_e5cabedd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[3]));
  AL_DFF_X al_ef3cfca0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[4]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[4]));
  AL_DFF_X al_9bfdb1da (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[5]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[5]));
  AL_DFF_X al_c25b66f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[6]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[6]));
  AL_DFF_X al_1be8e623 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b084da19[7]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5305cb61[7]));
  AL_DFF_X al_d1d228e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_df9b9d5b[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_e31e36f5[2]));
  AL_DFF_X al_b19106f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5743d58d[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_18d64456[0]));
  AL_DFF_X al_95b0bb1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5743d58d[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_18d64456[1]));
  AL_DFF_X al_2c0c4272 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5743d58d[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_18d64456[2]));
  AL_DFF_X al_107e7a90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5743d58d[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_18d64456[3]));
  AL_DFF_X al_1f47836d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5743d58d[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_18d64456[4]));
  AL_DFF_X al_618b1cd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5743d58d[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_18d64456[5]));
  AL_DFF_X al_82067f70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5743d58d[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_18d64456[6]));
  AL_DFF_X al_734c4999 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5743d58d[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_18d64456[7]));
  AL_DFF_X al_4cf0f6df (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[0]),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_6a6d2547[0]));
  AL_DFF_X al_8d09b7e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[1]),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_6a6d2547[1]));
  AL_DFF_X al_73f14769 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[2]),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_6a6d2547[2]));
  AL_DFF_X al_2534c1dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[3]),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_6a6d2547[3]));
  AL_DFF_X al_5144157b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[4]),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_6a6d2547[4]));
  AL_DFF_X al_f6832475 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[5]),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_6a6d2547[5]));
  AL_DFF_X al_e84cd853 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[6]),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_6a6d2547[6]));
  AL_DFF_X al_9d053fa5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[7]),
    .en(al_86ce862e),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_6a6d2547[7]));
  AL_DFF_X al_a03980f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e49f5b3[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ac23457[0]));
  AL_DFF_X al_89c380c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e49f5b3[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ac23457[1]));
  AL_DFF_X al_a193a498 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e49f5b3[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ac23457[2]));
  AL_DFF_X al_ab13b034 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e49f5b3[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ac23457[3]));
  AL_DFF_X al_679280f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e49f5b3[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ac23457[4]));
  AL_DFF_X al_2f9385d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e49f5b3[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ac23457[5]));
  AL_DFF_X al_32e320ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e49f5b3[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ac23457[6]));
  AL_DFF_X al_3fe7ba02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e49f5b3[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ac23457[7]));
  AL_DFF_X al_cde39bd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_30c5253d[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_1fc5093b[0]));
  AL_DFF_X al_89fbd83e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_21330e1d[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_1fc5093b[1]));
  AL_DFF_X al_caeec10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_21330e1d[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_1fc5093b[2]));
  AL_DFF_X al_7ef7d9b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_21330e1d[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_1fc5093b[3]));
  AL_DFF_X al_753e2645 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9bde74c4[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ab98f26[0]));
  AL_DFF_X al_f80afa80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9bde74c4[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_3ab98f26[1]));
  AL_DFF_X al_6025ca9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e44f12e[8]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ce55a07[8]));
  AL_DFF_X al_39f97cad (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e44f12e[9]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ce55a07[9]));
  AL_DFF_X al_998ddb6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e44f12e[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ce55a07[0]));
  AL_DFF_X al_c774d8ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e44f12e[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ce55a07[1]));
  AL_DFF_X al_93855ced (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e44f12e[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ce55a07[2]));
  AL_DFF_X al_b8df0bf8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e44f12e[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ce55a07[3]));
  AL_DFF_X al_8c7794dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e44f12e[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ce55a07[4]));
  AL_DFF_X al_4a93ad3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e44f12e[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ce55a07[5]));
  AL_DFF_X al_c2fd2da1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e44f12e[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ce55a07[6]));
  AL_DFF_X al_76fd25e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2e44f12e[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_3ce55a07[7]));
  AL_DFF_X al_d5f9f3bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[8]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_332a045d[8]));
  AL_DFF_X al_bce43c8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[9]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_332a045d[9]));
  AL_DFF_X al_29ff96c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[10]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_332a045d[10]));
  AL_DFF_X al_677dfae2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[11]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_332a045d[11]));
  AL_DFF_X al_5b28a33a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[12]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_332a045d[12]));
  AL_DFF_X al_5996bc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[13]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_332a045d[13]));
  AL_DFF_X al_94987a95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[14]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_332a045d[14]));
  AL_DFF_X al_a5a01961 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[15]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_332a045d[15]));
  AL_DFF_X al_5ab5241 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[16]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_332a045d[16]));
  AL_DFF_X al_5caec66a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[17]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_332a045d[17]));
  AL_DFF_X al_4f0ebfb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_332a045d[0]));
  AL_DFF_X al_ab3d2523 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[18]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_332a045d[18]));
  AL_DFF_X al_fd3a9fc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_332a045d[1]));
  AL_DFF_X al_5f647320 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_332a045d[2]));
  AL_DFF_X al_d95ec3f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_332a045d[3]));
  AL_DFF_X al_8dfe7e5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[4]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_332a045d[4]));
  AL_DFF_X al_ffb2e1cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[5]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_332a045d[5]));
  AL_DFF_X al_495146f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[6]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_332a045d[6]));
  AL_DFF_X al_bacde012 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dbdaab6[7]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_332a045d[7]));
  AL_DFF_X al_b428956c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ea27c82[0]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[8]));
  AL_DFF_X al_f709cde0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ea27c82[1]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[9]));
  AL_DFF_X al_174d4be8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ea27c82[2]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[10]));
  AL_DFF_X al_8cf7094f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ea27c82[3]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[11]));
  AL_DFF_X al_3d6641c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ea27c82[4]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[12]));
  AL_DFF_X al_1337b12e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ea27c82[5]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[13]));
  AL_DFF_X al_7e8d2138 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ea27c82[6]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[14]));
  AL_DFF_X al_8cb76138 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2ea27c82[7]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[15]));
  AL_DFF_X al_12e2c83e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f5fe9553[0]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[0]));
  AL_DFF_X al_b6e12b67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f5fe9553[1]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[1]));
  AL_DFF_X al_2682be7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f5fe9553[2]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[2]));
  AL_DFF_X al_c5acab47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f5fe9553[3]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[3]));
  AL_DFF_X al_a3192488 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f5fe9553[4]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[4]));
  AL_DFF_X al_b920f51a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f5fe9553[5]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[5]));
  AL_DFF_X al_15536524 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f5fe9553[6]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[6]));
  AL_DFF_X al_dcaaec86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f5fe9553[7]),
    .en(al_221dcc8d),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_eb2b30c3[7]));
  AL_DFF_X al_14d6f1de (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[8]));
  AL_DFF_X al_e5ea4825 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[8]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[9]));
  AL_DFF_X al_855239da (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[9]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[10]));
  AL_DFF_X al_f7d7c53c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[10]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[11]));
  AL_DFF_X al_52d0c4b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[11]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[12]));
  AL_DFF_X al_167424dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[12]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[13]));
  AL_DFF_X al_df6a6641 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd9f7a57),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[1]));
  AL_DFF_X al_c1af439f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[2]));
  AL_DFF_X al_4fac72cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[3]));
  AL_DFF_X al_4e52adce (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[4]));
  AL_DFF_X al_5f7c8a03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[5]));
  AL_DFF_X al_6cf92cc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[6]));
  AL_DFF_X al_92eabd5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cb8cffb4[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_cb8cffb4[7]));
  AL_DFF_X al_20bb31cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cf2a0a44[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_2a1554ab[0]));
  AL_DFF_X al_f9fa49b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cf2a0a44[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_2a1554ab[1]));
  AL_DFF_X al_1a569884 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cf2a0a44[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_2a1554ab[2]));
  AL_DFF_X al_4f34ba78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[7]));
  AL_DFF_X al_515f49f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[8]));
  AL_DFF_X al_86a1ac43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[9]));
  AL_DFF_X al_ac3bf91c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[10]));
  AL_DFF_X al_353e0163 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[11]));
  AL_DFF_X al_f23f5ebb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[8]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[12]));
  AL_DFF_X al_1343c5d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[9]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[13]));
  AL_DFF_X al_5bd5243b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[10]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[14]));
  AL_DFF_X al_e0ccf5dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[11]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[15]));
  AL_DFF_X al_786b323a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[12]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[16]));
  AL_DFF_X al_c90c2c76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_78612548),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[0]));
  AL_DFF_X al_6fbd454e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[13]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[17]));
  AL_DFF_X al_9962785f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_58e1cc88),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[19]));
  AL_DFF_X al_8d174d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ef80f5cf),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[21]));
  AL_DFF_X al_d680ffce (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_84db8eae),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[22]));
  AL_DFF_X al_9ad40604 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5dda436f),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[23]));
  AL_DFF_X al_d443dad3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d8c8c74d),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[28]));
  AL_DFF_X al_b64e6b2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1fc5093b[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[24]));
  AL_DFF_X al_e3727233 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1fc5093b[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[25]));
  AL_DFF_X al_7b2749a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1fc5093b[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[26]));
  AL_DFF_X al_e4084d2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3e1dba29),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[1]));
  AL_DFF_X al_d3d004b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1fc5093b[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[27]));
  AL_DFF_X al_1d1cbdcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_71ed2e0a),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[2]));
  AL_DFF_X al_b49346ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2c24255b),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[20]));
  AL_DFF_X al_a9a809e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_862844a1),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[18]));
  AL_DFF_X al_e79f860e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[4]));
  AL_DFF_X al_c99f8c5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[5]));
  AL_DFF_X al_38a9f8d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d28bc9[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(tx_status_vector[6]));
  AL_DFF_X al_2852fd1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_bd8e6c56),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_931288d8[0]));
  AL_DFF_X al_e11381ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_931288d8[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_931288d8[1]));
  AL_DFF_X al_1298d30d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[8]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[8]));
  AL_DFF_X al_beaf86cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[9]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[9]));
  AL_DFF_X al_5db7173c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[10]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[10]));
  AL_DFF_X al_ce19c95a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[11]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[11]));
  AL_DFF_X al_4fb169e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[12]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[12]));
  AL_DFF_X al_90bb2d01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[13]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[13]));
  AL_DFF_X al_63878caf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[0]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[0]));
  AL_DFF_X al_3dad5120 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[1]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[1]));
  AL_DFF_X al_995c3b79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[2]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[2]));
  AL_DFF_X al_8baab1a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[0]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[0]));
  AL_DFF_X al_95cfcf3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[3]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[3]));
  AL_DFF_X al_178e167c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[4]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[4]));
  AL_DFF_X al_f01dff1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[5]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[5]));
  AL_DFF_X al_8c05ba88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[6]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[6]));
  AL_DFF_X al_93f16cba (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[7]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[7]));
  AL_DFF_X al_737b6e94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[8]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[8]));
  AL_DFF_X al_8b42d7f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[9]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[9]));
  AL_DFF_X al_b4dd0624 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[10]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[10]));
  AL_DFF_X al_2a6bee8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[11]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[11]));
  AL_DFF_X al_1267d601 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[12]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[12]));
  AL_DFF_X al_1a19fd61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[1]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[1]));
  AL_DFF_X al_63682bca (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17c3d18e[13]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_e29488b2[13]));
  AL_DFF_X al_2428fb6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[0]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[0]));
  AL_DFF_X al_bad1c056 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[1]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[1]));
  AL_DFF_X al_2203d866 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[2]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[2]));
  AL_DFF_X al_e98b9ecc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[3]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[3]));
  AL_DFF_X al_1bf65fa2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[4]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[4]));
  AL_DFF_X al_f0b82eb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[5]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[5]));
  AL_DFF_X al_511d4fc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[6]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[6]));
  AL_DFF_X al_9ba0a89a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[7]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[7]));
  AL_DFF_X al_97aa64ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[2]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[2]));
  AL_DFF_X al_caaae434 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[8]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[8]));
  AL_DFF_X al_eb72db62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[9]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[9]));
  AL_DFF_X al_ccf4b7a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[10]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[10]));
  AL_DFF_X al_37a7e894 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[11]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[11]));
  AL_DFF_X al_a338246d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[12]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[12]));
  AL_DFF_X al_b5cf9bee (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[13]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[13]));
  AL_DFF_X al_c20d2201 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5305cb61[14]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_618d6d02[14]));
  AL_DFF_X al_98f0f0e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[3]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[3]));
  AL_DFF_X al_b847a06c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[4]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[4]));
  AL_DFF_X al_15bd4063 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[5]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[5]));
  AL_DFF_X al_4e3f02e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[6]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[6]));
  AL_DFF_X al_de9a2878 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e29488b2[7]),
    .en(al_5ce3a1c4),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_1a83737a[7]));
  AL_DFF_X al_94c55453 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aea1aa30[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_321109d3[0]));
  AL_DFF_X al_89def02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aea1aa30[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_321109d3[1]));
  AL_DFF_X al_7fe25b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4228c99a[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2ea27c82[0]));
  AL_DFF_X al_9b9c57b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4228c99a[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2ea27c82[1]));
  AL_DFF_X al_ed9f212d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4228c99a[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2ea27c82[2]));
  AL_DFF_X al_c39a10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4228c99a[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2ea27c82[3]));
  AL_DFF_X al_4b14f47c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4228c99a[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2ea27c82[4]));
  AL_DFF_X al_9ac7ca51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4228c99a[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2ea27c82[5]));
  AL_DFF_X al_18f1c164 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4228c99a[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2ea27c82[6]));
  AL_DFF_X al_8d6070d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4228c99a[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2ea27c82[7]));
  AL_DFF_X al_dc4de314 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8b969422[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f5fe9553[0]));
  AL_DFF_X al_b17b232a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d275691c[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f5fe9553[1]));
  AL_DFF_X al_92f5c9e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8b969422[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f5fe9553[2]));
  AL_DFF_X al_d73afb50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d275691c[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f5fe9553[3]));
  AL_DFF_X al_1b9d33ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8b969422[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f5fe9553[4]));
  AL_DFF_X al_22762e61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d275691c[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f5fe9553[5]));
  AL_DFF_X al_c0daca80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8b969422[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f5fe9553[6]));
  AL_DFF_X al_aadbd31e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d275691c[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_f5fe9553[7]));
  AL_DFF_X al_b82b400 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_da791a9b[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_31841a5b[0]));
  AL_DFF_X al_101ea05a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_da791a9b[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_31841a5b[1]));
  AL_DFF_X al_65e3542f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_da791a9b[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_31841a5b[2]));
  AL_DFF_X al_e42a5548 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_da791a9b[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_31841a5b[3]));
  AL_DFF_X al_a02cb997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_da791a9b[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_31841a5b[4]));
  AL_DFF_X al_b2d325e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_da791a9b[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_31841a5b[5]));
  AL_DFF_X al_35863ea3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_da791a9b[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_31841a5b[6]));
  AL_DFF_X al_49347c53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_da791a9b[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_31841a5b[7]));
  AL_DFF_X al_925a690e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_47ab7609[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d567b233[0]));
  AL_DFF_X al_588441a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_47ab7609[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d567b233[1]));
  AL_DFF_X al_304629b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_47ab7609[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d567b233[2]));
  AL_DFF_X al_2f77f9bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_47ab7609[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d567b233[3]));
  AL_DFF_X al_b9463117 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_47ab7609[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d567b233[4]));
  AL_DFF_X al_bbbc2e1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_47ab7609[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d567b233[5]));
  AL_DFF_X al_1e4d90f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_47ab7609[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d567b233[6]));
  AL_DFF_X al_749361f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_47ab7609[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_d567b233[7]));
  AL_DFF_X al_d6d23b8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d1fcb50b[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2453f186[0]));
  AL_DFF_X al_f2d6ffb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d1fcb50b[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2453f186[1]));
  AL_DFF_X al_be9c19ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d1fcb50b[2]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2453f186[2]));
  AL_DFF_X al_498cf1fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d1fcb50b[3]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2453f186[3]));
  AL_DFF_X al_46ca019c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d1fcb50b[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2453f186[4]));
  AL_DFF_X al_9308030 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d1fcb50b[5]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2453f186[5]));
  AL_DFF_X al_bfe28f15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d1fcb50b[6]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2453f186[6]));
  AL_DFF_X al_37590f75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d1fcb50b[7]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_2453f186[7]));
  AL_DFF_X al_f76f39c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[8]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_59a6ee8e[8]));
  AL_DFF_X al_764a46be (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[9]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_59a6ee8e[9]));
  AL_DFF_X al_d2e503f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[10]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_59a6ee8e[10]));
  AL_DFF_X al_23a11fec (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[11]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_59a6ee8e[11]));
  AL_DFF_X al_505da386 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[12]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_59a6ee8e[12]));
  AL_DFF_X al_eacbad69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[13]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_59a6ee8e[13]));
  AL_DFF_X al_9837e438 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[14]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_59a6ee8e[14]));
  AL_DFF_X al_1729e58f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[0]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_59a6ee8e[0]));
  AL_DFF_X al_bab7f2e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[1]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_59a6ee8e[1]));
  AL_DFF_X al_288baa8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_59a6ee8e[2]));
  AL_DFF_X al_f67ac2e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_59a6ee8e[3]));
  AL_DFF_X al_55d7a47b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[4]),
    .en(tx_clk_en),
    .sr(al_2dbca608),
    .ss(1'b0),
    .q(al_59a6ee8e[4]));
  AL_DFF_X al_9c764033 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[5]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_59a6ee8e[5]));
  AL_DFF_X al_a72559ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[6]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_59a6ee8e[6]));
  AL_DFF_X al_ff2631f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_49200bab[7]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_2dbca608),
    .q(al_59a6ee8e[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_74940e9 (
    .a(1'b0),
    .o({al_396e35f3,open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a0d00405 (
    .a(al_59a6ee8e[0]),
    .b(1'b1),
    .c(al_396e35f3),
    .o({al_c34e4fd4,al_83a6bf62[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3fc0e4e6 (
    .a(al_59a6ee8e[1]),
    .b(1'b0),
    .c(al_c34e4fd4),
    .o({al_57958b12,al_83a6bf62[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bf16ff0 (
    .a(al_59a6ee8e[2]),
    .b(1'b0),
    .c(al_57958b12),
    .o({al_3d6f4ec0,al_83a6bf62[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9d7b3ab6 (
    .a(al_59a6ee8e[3]),
    .b(1'b0),
    .c(al_3d6f4ec0),
    .o({al_7dd043ee,al_83a6bf62[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d30fab97 (
    .a(al_59a6ee8e[4]),
    .b(1'b0),
    .c(al_7dd043ee),
    .o({al_3226aea6,al_83a6bf62[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_79474cb0 (
    .a(al_59a6ee8e[5]),
    .b(1'b0),
    .c(al_3226aea6),
    .o({al_54e1a5bd,al_83a6bf62[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e44fa40f (
    .a(al_59a6ee8e[6]),
    .b(1'b0),
    .c(al_54e1a5bd),
    .o({al_9d8455d9,al_83a6bf62[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3a73d89b (
    .a(al_59a6ee8e[7]),
    .b(1'b0),
    .c(al_9d8455d9),
    .o({al_7a415511,al_83a6bf62[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fdbb04f3 (
    .a(al_59a6ee8e[8]),
    .b(1'b0),
    .c(al_7a415511),
    .o({al_26f9894f,al_83a6bf62[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27af8957 (
    .a(al_59a6ee8e[9]),
    .b(1'b0),
    .c(al_26f9894f),
    .o({al_ef281c2d,al_83a6bf62[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3b56d333 (
    .a(al_59a6ee8e[10]),
    .b(1'b0),
    .c(al_ef281c2d),
    .o({al_1db814d4,al_83a6bf62[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_966b475 (
    .a(al_59a6ee8e[11]),
    .b(1'b0),
    .c(al_1db814d4),
    .o({al_525a0f14,al_83a6bf62[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ce043e91 (
    .a(al_59a6ee8e[12]),
    .b(1'b0),
    .c(al_525a0f14),
    .o({al_3829c8d6,al_83a6bf62[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5b8e7393 (
    .a(al_59a6ee8e[13]),
    .b(1'b0),
    .c(al_3829c8d6),
    .o({al_c5560662,al_83a6bf62[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fdc09786 (
    .a(al_59a6ee8e[14]),
    .b(1'b0),
    .c(al_c5560662),
    .o({open_n19,al_83a6bf62[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_6d6b7eef (
    .a(1'b0),
    .o({al_26c32275,open_n22}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_32e10c9c (
    .a(al_332a045d[0]),
    .b(1'b1),
    .c(al_26c32275),
    .o({al_df53a2ee,al_cc156ef4[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_619b91f9 (
    .a(al_332a045d[1]),
    .b(1'b0),
    .c(al_df53a2ee),
    .o({al_a0dade4c,al_cc156ef4[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3b1f6115 (
    .a(al_332a045d[2]),
    .b(1'b0),
    .c(al_a0dade4c),
    .o({al_eb84a31d,al_cc156ef4[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_33d484ec (
    .a(al_332a045d[3]),
    .b(1'b0),
    .c(al_eb84a31d),
    .o({al_fe26d7bb,al_cc156ef4[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_67fc7040 (
    .a(al_332a045d[4]),
    .b(1'b0),
    .c(al_fe26d7bb),
    .o({al_7a228cbe,al_cc156ef4[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f0d285ba (
    .a(al_332a045d[5]),
    .b(1'b0),
    .c(al_7a228cbe),
    .o({al_be8ce4c3,al_cc156ef4[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8ab7dc2b (
    .a(al_332a045d[6]),
    .b(1'b0),
    .c(al_be8ce4c3),
    .o({al_bdda766f,al_cc156ef4[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7493dfd8 (
    .a(al_332a045d[7]),
    .b(1'b0),
    .c(al_bdda766f),
    .o({al_16346f67,al_cc156ef4[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b5725fc2 (
    .a(al_332a045d[8]),
    .b(1'b0),
    .c(al_16346f67),
    .o({al_90aba52e,al_cc156ef4[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_120c792a (
    .a(al_332a045d[9]),
    .b(1'b0),
    .c(al_90aba52e),
    .o({al_b4b4f932,al_cc156ef4[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f95d890c (
    .a(al_332a045d[10]),
    .b(1'b0),
    .c(al_b4b4f932),
    .o({al_39bec123,al_cc156ef4[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1c2d7c85 (
    .a(al_332a045d[11]),
    .b(1'b0),
    .c(al_39bec123),
    .o({al_6819cc15,al_cc156ef4[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_87554fe3 (
    .a(al_332a045d[12]),
    .b(1'b0),
    .c(al_6819cc15),
    .o({al_22cdf2f,al_cc156ef4[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_57d8ffa5 (
    .a(al_332a045d[13]),
    .b(1'b0),
    .c(al_22cdf2f),
    .o({al_1c995ac6,al_cc156ef4[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_48118d4b (
    .a(al_332a045d[14]),
    .b(1'b0),
    .c(al_1c995ac6),
    .o({al_2ef83128,al_cc156ef4[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d1b6b63c (
    .a(al_332a045d[15]),
    .b(1'b0),
    .c(al_2ef83128),
    .o({al_2cadd0ad,al_cc156ef4[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_82e8dca3 (
    .a(al_332a045d[16]),
    .b(1'b0),
    .c(al_2cadd0ad),
    .o({al_facb0130,al_cc156ef4[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6a6c9b71 (
    .a(al_332a045d[17]),
    .b(1'b0),
    .c(al_facb0130),
    .o({al_3bd7786d,al_cc156ef4[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5122109 (
    .a(al_332a045d[18]),
    .b(1'b0),
    .c(al_3bd7786d),
    .o({open_n23,al_cc156ef4[18]}));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_cabb9e07 (
    .a(al_7dd23876),
    .b(al_32c99495[3]),
    .o(al_b0d5abbb));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_270baa34 (
    .a(al_c4d87e5a),
    .b(al_859e5564),
    .c(al_7f22fda0),
    .d(al_4e2b6f95),
    .e(al_96662c62),
    .f(al_182d4638),
    .o(al_bd7f0fdb));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(C)*~(D)*~((~E*B))+~(A)*C*~(D)*~((~E*B))+A*C*~(D)*~((~E*B))+~(A)*~(C)*D*~((~E*B))+A*~(C)*D*~((~E*B))+~(A)*C*D*~((~E*B))+A*C*D*~((~E*B))+~(A)*~(C)*~(D)*(~E*B)+~(A)*C*~(D)*(~E*B)+A*C*~(D)*(~E*B)+~(A)*~(C)*D*(~E*B)+A*~(C)*D*(~E*B))"),
    .INIT(32'hfff53ff5))
    al_f64ea378 (
    .a(al_9e8adc84),
    .b(al_bd7f0fdb),
    .c(al_7f29f8c[1]),
    .d(al_7f29f8c[2]),
    .e(al_8213bac0),
    .o(al_1bd7127));
  AL_MAP_LUT5 #(
    .EQN("(A*B*~(C)*~((E*D))+~(A)*B*C*~((E*D))+A*B*C*~((E*D))+A*~(B)*~(C)*(E*D)+A*B*~(C)*(E*D)+~(A)*B*C*(E*D)+A*B*C*(E*D))"),
    .INIT(32'hcac8c8c8))
    al_42765699 (
    .a(al_1bd7127),
    .b(al_a6104abc),
    .c(al_7f29f8c[0]),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .o(al_271d4011));
  AL_DFF_X al_301cd991 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_271d4011),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_a6104abc));
  AL_MAP_LUT6 #(
    .EQN("(E*D*C*B*~(~F*~A))"),
    .INIT(64'hc000000080000000))
    al_ccef61a0 (
    .a(al_9e8adc84),
    .b(al_8f689368),
    .c(al_583c216b[1]),
    .d(al_583c216b[3]),
    .e(al_583c216b[5]),
    .f(al_c4d87e5a),
    .o(al_56237b7));
  AL_DFF_X al_2b2690a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_56237b7),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_c4d87e5a));
  AL_MAP_LUT6 #(
    .EQN("(~A*(C*~(B)*~((F*E*~D))+C*B*~((F*E*~D))+~(C)*B*(F*E*~D)+C*B*(F*E*~D)))"),
    .INIT(64'h5044505050505050))
    al_f4ed8f6c (
    .a(al_9e8adc84),
    .b(al_c4d87e5a),
    .c(al_bf03de15),
    .d(al_7f29f8c[0]),
    .e(al_7f29f8c[1]),
    .f(al_7f29f8c[2]),
    .o(al_af6ff858));
  AL_DFF_X al_c7ec8b34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_af6ff858),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_bf03de15));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~((~(~E*~D)*~C))+~(A)*~(B)*(~(~E*~D)*~C)+A*~(B)*(~(~E*~D)*~C)+A*B*(~(~E*~D)*~C))"),
    .INIT(32'h2b2b2b22))
    al_f23a267c (
    .a(al_d50b6ef8),
    .b(al_5f463be1),
    .c(al_7f29f8c[0]),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .o(al_abfa408b[0]));
  AL_MAP_LUT4 #(
    .EQN("((D@C)*~(B@A))"),
    .INIT(16'h0990))
    al_64c681b2 (
    .a(al_d50b6ef8),
    .b(al_5f463be1),
    .c(al_7f29f8c[0]),
    .d(al_7f29f8c[1]),
    .o(al_abfa408b[1]));
  AL_MAP_LUT5 #(
    .EQN("((E@(D*C))*~(B@A))"),
    .INIT(32'h09999000))
    al_5f4aea80 (
    .a(al_d50b6ef8),
    .b(al_5f463be1),
    .c(al_7f29f8c[0]),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .o(al_abfa408b[2]));
  AL_DFF_X al_e7775b64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d50b6ef8),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_5f463be1));
  AL_DFF_0 al_7c55335b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4c1d19df),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a2b89f7[0]));
  AL_DFF_0 al_187bd6a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6a2b89f7[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a2b89f7[1]));
  AL_DFF_0 al_a9b48996 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6a2b89f7[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a2b89f7[2]));
  AL_DFF_0 al_83ad1752 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6a2b89f7[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a2b89f7[3]));
  AL_DFF_0 al_1caa9dce (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_acd7ad28),
    .en(1'b1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_a927014c));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    al_83e461bd (
    .a(al_eb5eeaf9[4]),
    .b(al_eb5eeaf9[5]),
    .c(al_eb5eeaf9[6]),
    .d(al_eb5eeaf9[7]),
    .o(al_acd7ad28));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_cdf09aff (
    .a(al_5ffd8cb3[6]),
    .b(al_5ffd8cb3[14]),
    .c(al_5ffd8cb3[22]),
    .d(al_5ffd8cb3[30]),
    .e(al_7f29f8c[0]),
    .f(al_7f29f8c[1]),
    .o(al_8a20aaa));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(32'h00ca0000))
    al_d7265536 (
    .a(al_5ffd8cb3[33]),
    .b(al_5ffd8cb3[41]),
    .c(al_7f29f8c[0]),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .o(al_4d4393c7));
  AL_MAP_LUT5 #(
    .EQN("(C*~(B*A*~(E*D)))"),
    .INIT(32'hf0707070))
    al_2cd70ce7 (
    .a(al_dd43c64f),
    .b(al_d83e61fb),
    .c(al_5ffd8cb3[1]),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .o(al_d0651bd8));
  AL_MAP_LUT6 #(
    .EQN("(E@(~C*~(D*~(~B*~(~F*~A)))))"),
    .INIT(64'hfcf0030ffdf0020f))
    al_d148cecb (
    .a(al_a2fcb15d),
    .b(al_4d4393c7),
    .c(al_d0651bd8),
    .d(al_d50b6ef8),
    .e(al_583c216b[1]),
    .f(al_7f29f8c[2]),
    .o(al_b77a14d7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_3499771b (
    .a(al_5ffd8cb3[2]),
    .b(al_5ffd8cb3[10]),
    .c(al_5ffd8cb3[18]),
    .d(al_5ffd8cb3[26]),
    .e(al_7f29f8c[0]),
    .f(al_7f29f8c[1]),
    .o(al_8744257b));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d90a872f (
    .a(al_5ffd8cb3[34]),
    .b(al_5ffd8cb3[42]),
    .c(al_7f29f8c[0]),
    .o(al_aa714f0f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00cfc05f505f50))
    al_6ef89ef1 (
    .a(al_8744257b),
    .b(al_aa714f0f),
    .c(al_d50b6ef8),
    .d(al_5ffd8cb3[2]),
    .e(al_7f29f8c[1]),
    .f(al_7f29f8c[2]),
    .o(al_d7778ec8[2]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_a1e7e36a (
    .a(al_5ffd8cb3[3]),
    .b(al_5ffd8cb3[11]),
    .c(al_5ffd8cb3[19]),
    .d(al_5ffd8cb3[27]),
    .e(al_7f29f8c[0]),
    .f(al_7f29f8c[1]),
    .o(al_ded15eae));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_38a210f3 (
    .a(al_5ffd8cb3[35]),
    .b(al_5ffd8cb3[43]),
    .c(al_7f29f8c[0]),
    .o(al_50654b35));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00cfc05f505f50))
    al_5452947b (
    .a(al_ded15eae),
    .b(al_50654b35),
    .c(al_d50b6ef8),
    .d(al_5ffd8cb3[3]),
    .e(al_7f29f8c[1]),
    .f(al_7f29f8c[2]),
    .o(al_d7778ec8[3]));
  AL_MAP_LUT6 #(
    .EQN("(B*~A*~(F@D)*~(E@C))"),
    .INIT(64'h4000040000400004))
    al_7883e281 (
    .a(al_637261f7),
    .b(al_b77a14d7),
    .c(al_d7778ec8[2]),
    .d(al_d7778ec8[3]),
    .e(al_583c216b[2]),
    .f(al_583c216b[3]),
    .o(al_137e8f12));
  AL_MAP_LUT6 #(
    .EQN("(~E*(A*~(B)*~(C)*D*~(F)+A*B*~(C)*D*~(F)+A*~(B)*C*D*~(F)+A*B*C*D*~(F)+~(A)*B*~(C)*~(D)*F+A*B*~(C)*~(D)*F+~(A)*B*C*~(D)*F+A*B*C*~(D)*F+~(A)*~(B)*C*D*F+A*~(B)*C*D*F+~(A)*B*C*D*F+A*B*C*D*F))"),
    .INIT(64'h0000f0cc0000aa00))
    al_4baf3fc8 (
    .a(al_5ffd8cb3[13]),
    .b(al_5ffd8cb3[37]),
    .c(al_5ffd8cb3[45]),
    .d(al_7f29f8c[0]),
    .e(al_7f29f8c[1]),
    .f(al_7f29f8c[2]),
    .o(al_2408cdae));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F)"),
    .INIT(64'h5555ffff0f33ff55))
    al_d787ab6b (
    .a(al_5ffd8cb3[5]),
    .b(al_5ffd8cb3[21]),
    .c(al_5ffd8cb3[29]),
    .d(al_7f29f8c[0]),
    .e(al_7f29f8c[1]),
    .f(al_7f29f8c[2]),
    .o(al_a63c88b4));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(32'h00350000))
    al_8b87cfe7 (
    .a(al_5ffd8cb3[38]),
    .b(al_5ffd8cb3[46]),
    .c(al_7f29f8c[0]),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .o(al_b4bb4546));
  AL_MAP_LUT5 #(
    .EQN("(D@~(~E*~((B*~A))*~(C)+~E*(B*~A)*~(C)+~(~E)*(B*~A)*C+~E*(B*~A)*C))"),
    .INIT(32'h40bf4fb0))
    al_34952446 (
    .a(al_2408cdae),
    .b(al_a63c88b4),
    .c(al_d50b6ef8),
    .d(al_583c216b[5]),
    .e(al_5ffd8cb3[5]),
    .o(al_cc7e8768));
  AL_MAP_LUT6 #(
    .EQN("(~E*(A*~(B)*~(C)*D*~(F)+A*B*~(C)*D*~(F)+A*~(B)*C*D*~(F)+A*B*C*D*~(F)+~(A)*B*~(C)*~(D)*F+A*B*~(C)*~(D)*F+~(A)*B*C*~(D)*F+A*B*C*~(D)*F+~(A)*~(B)*C*D*F+A*~(B)*C*D*F+~(A)*B*C*D*F+A*B*C*D*F))"),
    .INIT(64'h0000f0cc0000aa00))
    al_113da2ef (
    .a(al_5ffd8cb3[8]),
    .b(al_5ffd8cb3[32]),
    .c(al_5ffd8cb3[40]),
    .d(al_7f29f8c[0]),
    .e(al_7f29f8c[1]),
    .f(al_7f29f8c[2]),
    .o(al_83be6442));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+~(A)*B*C*D*E*F)"),
    .INIT(64'h5555ffff0f33ff55))
    al_b38ec0bb (
    .a(al_5ffd8cb3[0]),
    .b(al_5ffd8cb3[16]),
    .c(al_5ffd8cb3[24]),
    .d(al_7f29f8c[0]),
    .e(al_7f29f8c[1]),
    .f(al_7f29f8c[2]),
    .o(al_b0d20bea));
  AL_MAP_LUT5 #(
    .EQN("(D@~(~E*~((B*~A))*~(C)+~E*(B*~A)*~(C)+~(~E)*(B*~A)*C+~E*(B*~A)*C))"),
    .INIT(32'h40bf4fb0))
    al_d93def0c (
    .a(al_83be6442),
    .b(al_b0d20bea),
    .c(al_d50b6ef8),
    .d(al_583c216b[0]),
    .e(al_5ffd8cb3[0]),
    .o(al_76c6b29d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_63ac1f45 (
    .a(al_5ffd8cb3[4]),
    .b(al_5ffd8cb3[12]),
    .c(al_5ffd8cb3[20]),
    .d(al_5ffd8cb3[28]),
    .e(al_7f29f8c[0]),
    .f(al_7f29f8c[1]),
    .o(al_98c88117));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5e014f2f (
    .a(al_5ffd8cb3[36]),
    .b(al_5ffd8cb3[44]),
    .c(al_7f29f8c[0]),
    .o(al_554dd8ee));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00cfc05f505f50))
    al_934854c6 (
    .a(al_98c88117),
    .b(al_554dd8ee),
    .c(al_d50b6ef8),
    .d(al_5ffd8cb3[4]),
    .e(al_7f29f8c[1]),
    .f(al_7f29f8c[2]),
    .o(al_d7778ec8[4]));
  AL_MAP_LUT5 #(
    .EQN("(E*~B*~A*~(D@C))"),
    .INIT(32'h10010000))
    al_708b42bc (
    .a(al_cc7e8768),
    .b(al_76c6b29d),
    .c(al_d7778ec8[4]),
    .d(al_583c216b[4]),
    .e(al_859e5564),
    .o(al_4a2c328a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_1b819e78 (
    .a(al_5ffd8cb3[7]),
    .b(al_5ffd8cb3[15]),
    .c(al_5ffd8cb3[23]),
    .d(al_5ffd8cb3[31]),
    .e(al_7f29f8c[0]),
    .f(al_7f29f8c[1]),
    .o(al_ec1c3fd8));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h020e323ec2cef2fe))
    al_36f0876a (
    .a(al_ec1c3fd8),
    .b(al_d7f7aaa1),
    .c(al_c2044b3b),
    .d(al_5ffd8cb3[7]),
    .e(al_5ffd8cb3[39]),
    .f(al_5ffd8cb3[47]),
    .o(al_8c91da92));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_f8661e94 (
    .a(al_8c91da92),
    .b(al_d50b6ef8),
    .c(al_5ffd8cb3[7]),
    .o(al_d7778ec8[7]));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(B*A*~(E@C)))"),
    .INIT(32'hff80ff08))
    al_a7eb4917 (
    .a(al_137e8f12),
    .b(al_4a2c328a),
    .c(al_d7778ec8[7]),
    .d(al_dbd06164),
    .e(al_583c216b[7]),
    .o(al_772d3492));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(B*A*~(E*D)))"),
    .INIT(32'h0f070707))
    al_2990ee4f (
    .a(al_dd43c64f),
    .b(al_d83e61fb),
    .c(al_5ffd8cb3[6]),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .o(al_d2a71eb2));
  AL_MAP_LUT6 #(
    .EQN("(E@(~C*~(D*~(~B*~(~F*A)))))"),
    .INIT(64'hfcf0030ffef0010f))
    al_be458259 (
    .a(al_8a20aaa),
    .b(al_b4bb4546),
    .c(al_d2a71eb2),
    .d(al_d50b6ef8),
    .e(al_583c216b[6]),
    .f(al_7f29f8c[2]),
    .o(al_637261f7));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00ff0f0f33335555))
    al_b6ffa628 (
    .a(al_5ffd8cb3[1]),
    .b(al_5ffd8cb3[9]),
    .c(al_5ffd8cb3[17]),
    .d(al_5ffd8cb3[25]),
    .e(al_7f29f8c[0]),
    .f(al_7f29f8c[1]),
    .o(al_a2fcb15d));
  AL_DFF_X al_9af20628 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_772d3492),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_859e5564));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_e1013fdc (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_b7012aee[5]),
    .d(al_b7012aee[13]),
    .e(al_b7012aee[21]),
    .f(al_b7012aee[29]),
    .o(al_a808afa8));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*~(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))"),
    .INIT(32'h00102030))
    al_8d639704 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .d(al_b7012aee[38]),
    .e(al_b7012aee[46]),
    .o(al_8e9644e7));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(B*A*~(D*C)))"),
    .INIT(32'h0000f777))
    al_fef5dfb9 (
    .a(al_dd43c64f),
    .b(al_d83e61fb),
    .c(al_7f29f8c[1]),
    .d(al_7f29f8c[2]),
    .e(al_b7012aee[6]),
    .o(al_54a9598a));
  AL_MAP_LUT6 #(
    .EQN("(E@(~C*~(D*~(~B*~(~F*A)))))"),
    .INIT(64'hfcf0030ffef0010f))
    al_db700f82 (
    .a(al_3dc2993c),
    .b(al_8e9644e7),
    .c(al_54a9598a),
    .d(al_d50b6ef8),
    .e(al_583c216b[6]),
    .f(al_7f29f8c[2]),
    .o(al_aca9177e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_6c8f5c76 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_b7012aee[4]),
    .d(al_b7012aee[12]),
    .e(al_b7012aee[20]),
    .f(al_b7012aee[28]),
    .o(al_85f33b95));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_75e3f7bf (
    .a(al_7f29f8c[0]),
    .b(al_b7012aee[36]),
    .c(al_b7012aee[44]),
    .o(al_8345e39d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffcf5f5f00c05050))
    al_569d42ba (
    .a(al_85f33b95),
    .b(al_8345e39d),
    .c(al_d50b6ef8),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .f(al_b7012aee[4]),
    .o(al_d7778ec8[12]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_db7feb16 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_b7012aee[3]),
    .d(al_b7012aee[11]),
    .e(al_b7012aee[19]),
    .f(al_b7012aee[27]),
    .o(al_c03c1e89));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_33a93da8 (
    .a(al_7f29f8c[0]),
    .b(al_b7012aee[35]),
    .c(al_b7012aee[43]),
    .o(al_338c309a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffcf5f5f00c05050))
    al_acb7a96f (
    .a(al_c03c1e89),
    .b(al_338c309a),
    .c(al_d50b6ef8),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .f(al_b7012aee[3]),
    .o(al_d7778ec8[11]));
  AL_MAP_LUT6 #(
    .EQN("(~B*A*~(E@D)*~(F@C))"),
    .INIT(64'h2000002002000002))
    al_14ed05d0 (
    .a(al_999473bf),
    .b(al_aca9177e),
    .c(al_d7778ec8[12]),
    .d(al_d7778ec8[11]),
    .e(al_583c216b[3]),
    .f(al_583c216b[4]),
    .o(al_df93f3b6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_b9c15a9a (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_b7012aee[2]),
    .d(al_b7012aee[10]),
    .e(al_b7012aee[18]),
    .f(al_b7012aee[26]),
    .o(al_bc71b143));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bfc4fa21 (
    .a(al_7f29f8c[0]),
    .b(al_b7012aee[34]),
    .c(al_b7012aee[42]),
    .o(al_5f7aacbd));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffcf5f5f00c05050))
    al_2961f9e (
    .a(al_bc71b143),
    .b(al_5f7aacbd),
    .c(al_d50b6ef8),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .f(al_b7012aee[2]),
    .o(al_d7778ec8[10]));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))"),
    .INIT(32'h30201000))
    al_8dcda6d6 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .d(al_b7012aee[37]),
    .e(al_b7012aee[45]),
    .o(al_8a909a7e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_24104606 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_b7012aee[1]),
    .d(al_b7012aee[9]),
    .e(al_b7012aee[17]),
    .f(al_b7012aee[25]),
    .o(al_c6d8833c));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_34d04096 (
    .a(al_7f29f8c[0]),
    .b(al_b7012aee[33]),
    .c(al_b7012aee[41]),
    .o(al_51ce9e18));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffcf5f5f00c05050))
    al_d881d89e (
    .a(al_c6d8833c),
    .b(al_51ce9e18),
    .c(al_d50b6ef8),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .f(al_b7012aee[1]),
    .o(al_d7778ec8[9]));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    al_85db4fd (
    .a(al_d7778ec8[10]),
    .b(al_d7778ec8[9]),
    .c(al_583c216b[1]),
    .d(al_583c216b[2]),
    .o(al_abb85d9));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hcbcfdbdfebeffbff))
    al_4bdc3cef (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .d(al_b7012aee[23]),
    .e(al_b7012aee[39]),
    .f(al_b7012aee[47]),
    .o(al_4503fb38));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~((E*~(F)*~(C)+E*F*~(C)+~(E)*F*C+E*F*C))*~((~D*B))+~A*(E*~(F)*~(C)+E*F*~(C)+~(E)*F*C+E*F*C)*~((~D*B))+~(~A)*(E*~(F)*~(C)+E*F*~(C)+~(E)*F*C+E*F*C)*(~D*B)+~A*(E*~(F)*~(C)+E*F*~(C)+~(E)*F*C+E*F*C)*(~D*B))"),
    .INIT(64'haa22aa2eaae2aaee))
    al_3675370c (
    .a(al_4503fb38),
    .b(al_7f29f8c[0]),
    .c(al_7f29f8c[1]),
    .d(al_7f29f8c[2]),
    .e(al_b7012aee[15]),
    .f(al_b7012aee[31]),
    .o(al_8298897d));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*C*D)"),
    .INIT(16'h80af))
    al_cbafea8b (
    .a(al_8298897d),
    .b(al_34ca3fbe),
    .c(al_d50b6ef8),
    .d(al_b7012aee[7]),
    .o(al_56a26cfa));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfdb97531))
    al_9e6fa8ba (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_b7012aee[8]),
    .d(al_b7012aee[16]),
    .e(al_b7012aee[24]),
    .o(al_58887de));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~((~C*~(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))*~(D)+~A*(~C*~(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*~(D)+~(~A)*(~C*~(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*D+~A*(~C*~(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*D)"),
    .INIT(64'hffaafcaaf3aaf0aa))
    al_54e6febb (
    .a(al_58887de),
    .b(al_7f29f8c[0]),
    .c(al_7f29f8c[1]),
    .d(al_7f29f8c[2]),
    .e(al_b7012aee[32]),
    .f(al_b7012aee[40]),
    .o(al_9073553b));
  AL_MAP_LUT6 #(
    .EQN("(E*(D@(~(A)*~(B)*~(C)*~(F)+A*~(B)*~(C)*~(F)+~(A)*B*~(C)*~(F)+A*B*~(C)*~(F)+~(A)*~(B)*C*~(F)+A*~(B)*C*~(F)+~(A)*B*C*~(F)+~(A)*~(B)*C*F+~(A)*B*C*F)))"),
    .INIT(64'haf500000807f0000))
    al_8ccfe11a (
    .a(al_9073553b),
    .b(al_34ca3fbe),
    .c(al_d50b6ef8),
    .d(al_583c216b[0]),
    .e(al_7f22fda0),
    .f(al_b7012aee[0]),
    .o(al_d8b60780));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~(D*B*A*(F@C)))"),
    .INIT(64'hffff0800ffff8000))
    al_2ec06417 (
    .a(al_df93f3b6),
    .b(al_abb85d9),
    .c(al_56a26cfa),
    .d(al_d8b60780),
    .e(al_dbd06164),
    .f(al_583c216b[7]),
    .o(al_8af9f67c));
  AL_MAP_LUT5 #(
    .EQN("(E*~(B*A*~(D*C)))"),
    .INIT(32'hf7770000))
    al_32ade8d9 (
    .a(al_dd43c64f),
    .b(al_d83e61fb),
    .c(al_7f29f8c[1]),
    .d(al_7f29f8c[2]),
    .e(al_b7012aee[5]),
    .o(al_7a2b8846));
  AL_MAP_LUT6 #(
    .EQN("(E@(~C*~(D*~(~B*~(~F*~A)))))"),
    .INIT(64'hfcf0030ffdf0020f))
    al_7191a5eb (
    .a(al_a808afa8),
    .b(al_8a909a7e),
    .c(al_7a2b8846),
    .d(al_d50b6ef8),
    .e(al_583c216b[5]),
    .f(al_7f29f8c[2]),
    .o(al_999473bf));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_cef2695d (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_b7012aee[6]),
    .d(al_b7012aee[14]),
    .e(al_b7012aee[22]),
    .f(al_b7012aee[30]),
    .o(al_3dc2993c));
  AL_DFF_X al_a53375ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8af9f67c),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7f22fda0));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_156979f9 (
    .a(al_dd43c64f),
    .b(al_d83e61fb),
    .o(al_d50b6ef8));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_4d5beecf (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_f07b9ef6[0]),
    .d(al_f07b9ef6[8]),
    .e(al_f07b9ef6[16]),
    .f(al_f07b9ef6[24]),
    .o(al_4f0b110));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_620c5cf0 (
    .a(al_7f29f8c[0]),
    .b(al_f07b9ef6[32]),
    .c(al_f07b9ef6[40]),
    .o(al_d55c6f72));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F)"),
    .INIT(64'h0030a0a0ff3fafaf))
    al_5ca45a68 (
    .a(al_4f0b110),
    .b(al_d55c6f72),
    .c(al_d50b6ef8),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .f(al_f07b9ef6[0]),
    .o(al_ac502f3b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_de646b5a (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_f07b9ef6[1]),
    .d(al_f07b9ef6[9]),
    .e(al_f07b9ef6[17]),
    .f(al_f07b9ef6[25]),
    .o(al_b5cc7793));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_32f893b0 (
    .a(al_7f29f8c[0]),
    .b(al_f07b9ef6[33]),
    .c(al_f07b9ef6[41]),
    .o(al_37adc87c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffcf5f5f00c05050))
    al_7891969b (
    .a(al_b5cc7793),
    .b(al_37adc87c),
    .c(al_d50b6ef8),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .f(al_f07b9ef6[1]),
    .o(al_d7778ec8[17]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_3ad5a79a (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_f07b9ef6[5]),
    .d(al_f07b9ef6[13]),
    .e(al_f07b9ef6[21]),
    .f(al_f07b9ef6[29]),
    .o(al_503c8f93));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_e24ad424 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .o(al_d7f7aaa1));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_66f92c10 (
    .a(al_7f29f8c[0]),
    .b(al_f07b9ef6[37]),
    .c(al_f07b9ef6[45]),
    .o(al_c6b2b040));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hffcf5f5f00c05050))
    al_ef4f90c7 (
    .a(al_503c8f93),
    .b(al_c6b2b040),
    .c(al_d50b6ef8),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .f(al_f07b9ef6[5]),
    .o(al_d7778ec8[21]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*(D@A))"),
    .INIT(64'h4080102004080102))
    al_e6338937 (
    .a(al_ac502f3b),
    .b(al_d7778ec8[17]),
    .c(al_d7778ec8[21]),
    .d(al_583c216b[0]),
    .e(al_583c216b[1]),
    .f(al_583c216b[5]),
    .o(al_a81bacbe));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_e3c6ae8d (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .d(al_f07b9ef6[15]),
    .e(al_f07b9ef6[39]),
    .f(al_f07b9ef6[47]),
    .o(al_72c24a7e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h32f336f73afb3eff))
    al_81981f41 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .d(al_f07b9ef6[7]),
    .e(al_f07b9ef6[23]),
    .f(al_f07b9ef6[31]),
    .o(al_d67debd3));
  AL_MAP_LUT5 #(
    .EQN("(D@~(~E*~((B*~A))*~(C)+~E*(B*~A)*~(C)+~(~E)*(B*~A)*C+~E*(B*~A)*C))"),
    .INIT(32'h40bf4fb0))
    al_46deb39f (
    .a(al_72c24a7e),
    .b(al_d67debd3),
    .c(al_d50b6ef8),
    .d(al_583c216b[7]),
    .e(al_f07b9ef6[7]),
    .o(al_69d9a189));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_776cd1df (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .d(al_f07b9ef6[14]),
    .e(al_f07b9ef6[38]),
    .f(al_f07b9ef6[46]),
    .o(al_809052dd));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h32f336f73afb3eff))
    al_b32c056d (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .d(al_f07b9ef6[6]),
    .e(al_f07b9ef6[22]),
    .f(al_f07b9ef6[30]),
    .o(al_6be58e65));
  AL_MAP_LUT5 #(
    .EQN("(D@~(~E*~((B*~A))*~(C)+~E*(B*~A)*~(C)+~(~E)*(B*~A)*C+~E*(B*~A)*C))"),
    .INIT(32'h40bf4fb0))
    al_4f36741 (
    .a(al_809052dd),
    .b(al_6be58e65),
    .c(al_d50b6ef8),
    .d(al_583c216b[6]),
    .e(al_f07b9ef6[6]),
    .o(al_f5473a34));
  AL_MAP_LUT6 #(
    .EQN("(~C*(A*~(B)*D*~(E)*~(F)+~(A)*B*~(D)*E*~(F)+A*~(B)*D*E*~(F)+~(A)*B*D*E*~(F)+A*B*~(D)*~(E)*F+A*~(B)*D*~(E)*F+A*B*D*~(E)*F+~(A)*B*~(D)*E*F+A*B*~(D)*E*F+A*~(B)*D*E*F+~(A)*B*D*E*F+A*B*D*E*F))"),
    .INIT(64'h0e0c0a0806040200))
    al_4f787dee (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .d(al_f07b9ef6[11]),
    .e(al_f07b9ef6[19]),
    .f(al_f07b9ef6[27]),
    .o(al_95fe37a9));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))"),
    .INIT(32'h30201000))
    al_2373521 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .d(al_f07b9ef6[35]),
    .e(al_f07b9ef6[43]),
    .o(al_c8d005d));
  AL_MAP_LUT5 #(
    .EQN("(~((~B*~A))*~(C)*D*~(E)+~((~B*~A))*C*D*~(E)+~((~B*~A))*~(C)*~(D)*E+(~B*~A)*~(C)*~(D)*E+~((~B*~A))*C*~(D)*E+(~B*~A)*C*~(D)*E+~((~B*~A))*~(C)*D*E+(~B*~A)*~(C)*D*E+~((~B*~A))*C*D*E)"),
    .INIT(32'hefffee00))
    al_3443abb8 (
    .a(al_95fe37a9),
    .b(al_c8d005d),
    .c(al_34ca3fbe),
    .d(al_d50b6ef8),
    .e(al_f07b9ef6[3]),
    .o(al_d7778ec8[19]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_8fbbfd1c (
    .a(al_7f29f8c[1]),
    .b(al_7f29f8c[2]),
    .o(al_c2044b3b));
  AL_MAP_LUT5 #(
    .EQN("(E*~B*~A*~(D@C))"),
    .INIT(32'h10010000))
    al_5174946f (
    .a(al_69d9a189),
    .b(al_f5473a34),
    .c(al_d7778ec8[19]),
    .d(al_583c216b[3]),
    .e(al_4e2b6f95),
    .o(al_aacf80e2));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_430eb6ab (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_f07b9ef6[4]),
    .d(al_f07b9ef6[12]),
    .e(al_f07b9ef6[20]),
    .f(al_f07b9ef6[28]),
    .o(al_68eb24f8));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*~(C)*D*E*F)"),
    .INIT(64'h020e323ec2cef2fe))
    al_522f3078 (
    .a(al_68eb24f8),
    .b(al_d7f7aaa1),
    .c(al_c2044b3b),
    .d(al_f07b9ef6[4]),
    .e(al_f07b9ef6[36]),
    .f(al_f07b9ef6[44]),
    .o(al_a07f4463));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_ef92acf1 (
    .a(al_a07f4463),
    .b(al_d50b6ef8),
    .c(al_f07b9ef6[4]),
    .o(al_d7778ec8[20]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F)"),
    .INIT(64'h0123456789abcdef))
    al_34a36b89 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_f07b9ef6[2]),
    .d(al_f07b9ef6[10]),
    .e(al_f07b9ef6[18]),
    .f(al_f07b9ef6[26]),
    .o(al_78627e02));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8d762e51 (
    .a(al_7f29f8c[0]),
    .b(al_f07b9ef6[34]),
    .c(al_f07b9ef6[42]),
    .o(al_82d0eff2));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccfff5ffcc000500))
    al_6a23cfb5 (
    .a(al_78627e02),
    .b(al_82d0eff2),
    .c(al_d7f7aaa1),
    .d(al_d50b6ef8),
    .e(al_c2044b3b),
    .f(al_f07b9ef6[2]),
    .o(al_d7778ec8[18]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_c0cb02be (
    .a(al_d7778ec8[18]),
    .b(al_583c216b[2]),
    .o(al_bc4e38bd));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~(D*B*A*~(F@C)))"),
    .INIT(64'hffff8000ffff0800))
    al_d3192caa (
    .a(al_a81bacbe),
    .b(al_aacf80e2),
    .c(al_d7778ec8[20]),
    .d(al_bc4e38bd),
    .e(al_dbd06164),
    .f(al_583c216b[4]),
    .o(al_513305d5));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_cb96a5c2 (
    .a(al_d50b6ef8),
    .b(al_7f29f8c[0]),
    .c(al_7f29f8c[1]),
    .d(al_7f29f8c[2]),
    .o(al_dbd06164));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C)"),
    .INIT(8'h3e))
    al_9d827c08 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .o(al_34ca3fbe));
  AL_DFF_X al_18bee407 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_513305d5),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4e2b6f95));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_613c3352 (
    .a(s_axi_awvalid),
    .b(s_axi_wvalid),
    .c(s_axi_awready),
    .o(al_26874532));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_dbd15d21 (
    .a(al_26874532),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_c9ac0c17));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_efec4166 (
    .a(al_60c7c349[2]),
    .b(al_60c7c349[3]),
    .o(al_cc5f5ce9));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    al_1296e252 (
    .a(al_f931229[0]),
    .b(al_f931229[1]),
    .c(al_f931229[2]),
    .d(al_f931229[3]),
    .o(al_223a077f));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'h00800000))
    al_2b4a7984 (
    .a(al_c9ac0c17),
    .b(al_cc5f5ce9),
    .c(al_223a077f),
    .d(al_60c7c349[0]),
    .e(al_60c7c349[1]),
    .o(al_be4e813d));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_faf95db3 (
    .a(al_c9ac0c17),
    .b(al_cc5f5ce9),
    .c(al_223a077f),
    .d(al_60c7c349[0]),
    .e(al_60c7c349[1]),
    .o(al_d0f70766));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_e397f4f1 (
    .a(al_f931229[0]),
    .b(al_f931229[1]),
    .c(al_f931229[2]),
    .d(al_f931229[3]),
    .o(al_f44488cf));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'h00800000))
    al_e2729628 (
    .a(al_c9ac0c17),
    .b(al_cc5f5ce9),
    .c(al_f44488cf),
    .d(al_60c7c349[0]),
    .e(al_60c7c349[1]),
    .o(al_db3a7a8b));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_e337154b (
    .a(al_c9ac0c17),
    .b(al_cc5f5ce9),
    .c(al_f44488cf),
    .d(al_60c7c349[0]),
    .e(al_60c7c349[1]),
    .o(al_297252e3));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_2263b39d (
    .a(al_f931229[0]),
    .b(al_f931229[1]),
    .c(al_f931229[2]),
    .d(al_f931229[3]),
    .o(al_e7ad9386));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'h00800000))
    al_59ff2a2e (
    .a(al_c9ac0c17),
    .b(al_cc5f5ce9),
    .c(al_e7ad9386),
    .d(al_60c7c349[0]),
    .e(al_60c7c349[1]),
    .o(al_9e004fa1));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_7c72a36d (
    .a(al_c9ac0c17),
    .b(al_cc5f5ce9),
    .c(al_e7ad9386),
    .d(al_60c7c349[0]),
    .e(al_60c7c349[1]),
    .o(al_5a460c8d));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_eab61ffa (
    .a(al_d50b6ef8),
    .b(al_42381c95[0]),
    .c(al_b091d0de[8]),
    .o(al_e49fcd23[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_de78f9ad (
    .a(al_d50b6ef8),
    .b(al_42381c95[10]),
    .c(al_b091d0de[18]),
    .o(al_e49fcd23[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_622c4c4c (
    .a(al_d50b6ef8),
    .b(al_42381c95[11]),
    .c(al_b091d0de[19]),
    .o(al_e49fcd23[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c833474a (
    .a(al_d50b6ef8),
    .b(al_42381c95[12]),
    .c(al_b091d0de[20]),
    .o(al_e49fcd23[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4ce856d2 (
    .a(al_d50b6ef8),
    .b(al_42381c95[13]),
    .c(al_b091d0de[21]),
    .o(al_e49fcd23[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_da2c1525 (
    .a(al_d50b6ef8),
    .b(al_42381c95[14]),
    .c(al_b091d0de[22]),
    .o(al_e49fcd23[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_996d1e3d (
    .a(al_d50b6ef8),
    .b(al_42381c95[15]),
    .c(al_b091d0de[23]),
    .o(al_e49fcd23[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4499991b (
    .a(al_d50b6ef8),
    .b(al_42381c95[16]),
    .c(al_b091d0de[24]),
    .o(al_e49fcd23[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_eea38d18 (
    .a(al_d50b6ef8),
    .b(al_42381c95[17]),
    .c(al_b091d0de[25]),
    .o(al_e49fcd23[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2e8e9088 (
    .a(al_d50b6ef8),
    .b(al_42381c95[18]),
    .c(al_b091d0de[26]),
    .o(al_e49fcd23[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_91fa3f5e (
    .a(al_d50b6ef8),
    .b(al_42381c95[19]),
    .c(al_b091d0de[27]),
    .o(al_e49fcd23[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f03384e4 (
    .a(al_d50b6ef8),
    .b(al_42381c95[1]),
    .c(al_b091d0de[9]),
    .o(al_e49fcd23[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_202aad4b (
    .a(al_d50b6ef8),
    .b(al_42381c95[20]),
    .c(al_b091d0de[28]),
    .o(al_e49fcd23[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f0fac29a (
    .a(al_d50b6ef8),
    .b(al_42381c95[21]),
    .c(al_b091d0de[29]),
    .o(al_e49fcd23[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2329160 (
    .a(al_d50b6ef8),
    .b(al_42381c95[22]),
    .c(al_b091d0de[30]),
    .o(al_e49fcd23[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3c09b25c (
    .a(al_d50b6ef8),
    .b(al_42381c95[23]),
    .c(al_b091d0de[31]),
    .o(al_e49fcd23[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bc6bf736 (
    .a(al_d50b6ef8),
    .b(al_42381c95[24]),
    .c(al_b091d0de[32]),
    .o(al_e49fcd23[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bd64dab3 (
    .a(al_d50b6ef8),
    .b(al_42381c95[25]),
    .c(al_b091d0de[33]),
    .o(al_e49fcd23[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f09aae66 (
    .a(al_d50b6ef8),
    .b(al_42381c95[26]),
    .c(al_b091d0de[34]),
    .o(al_e49fcd23[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c4143918 (
    .a(al_d50b6ef8),
    .b(al_42381c95[27]),
    .c(al_b091d0de[35]),
    .o(al_e49fcd23[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_38d159fb (
    .a(al_d50b6ef8),
    .b(al_42381c95[28]),
    .c(al_b091d0de[36]),
    .o(al_e49fcd23[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_aed9ce95 (
    .a(al_d50b6ef8),
    .b(al_42381c95[29]),
    .c(al_b091d0de[37]),
    .o(al_e49fcd23[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_101fb691 (
    .a(al_d50b6ef8),
    .b(al_42381c95[2]),
    .c(al_b091d0de[10]),
    .o(al_e49fcd23[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b407cf78 (
    .a(al_d50b6ef8),
    .b(al_42381c95[30]),
    .c(al_b091d0de[38]),
    .o(al_e49fcd23[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7a721c2b (
    .a(al_d50b6ef8),
    .b(al_42381c95[31]),
    .c(al_b091d0de[39]),
    .o(al_e49fcd23[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_63509306 (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[0]),
    .c(al_b091d0de[40]),
    .o(al_e49fcd23[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_70492004 (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[1]),
    .c(al_b091d0de[41]),
    .o(al_e49fcd23[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c2ed2413 (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[2]),
    .c(al_b091d0de[42]),
    .o(al_e49fcd23[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_595f27eb (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[3]),
    .c(al_b091d0de[43]),
    .o(al_e49fcd23[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6ae15cd2 (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[4]),
    .c(al_b091d0de[44]),
    .o(al_e49fcd23[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d5cf1191 (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[5]),
    .c(al_b091d0de[45]),
    .o(al_e49fcd23[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9a6cdd2b (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[6]),
    .c(al_b091d0de[46]),
    .o(al_e49fcd23[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6681cac8 (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[7]),
    .c(al_b091d0de[47]),
    .o(al_e49fcd23[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2467bc53 (
    .a(al_d50b6ef8),
    .b(al_42381c95[3]),
    .c(al_b091d0de[11]),
    .o(al_e49fcd23[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_3987da4e (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[8]),
    .o(al_e49fcd23[40]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b8a66fba (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[9]),
    .o(al_e49fcd23[41]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_cedf74ea (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[10]),
    .o(al_e49fcd23[42]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_a1d24711 (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[11]),
    .o(al_e49fcd23[43]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_508b3201 (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[12]),
    .o(al_e49fcd23[44]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6e3ac8be (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[13]),
    .o(al_e49fcd23[45]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_25e1cbd (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[14]),
    .o(al_e49fcd23[46]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_139348a9 (
    .a(al_d50b6ef8),
    .b(al_a3c2ad2a[15]),
    .o(al_e49fcd23[47]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_89d8a7b (
    .a(al_d50b6ef8),
    .b(al_42381c95[4]),
    .c(al_b091d0de[12]),
    .o(al_e49fcd23[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2073c6a2 (
    .a(al_d50b6ef8),
    .b(al_42381c95[5]),
    .c(al_b091d0de[13]),
    .o(al_e49fcd23[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_181711c4 (
    .a(al_d50b6ef8),
    .b(al_42381c95[6]),
    .c(al_b091d0de[14]),
    .o(al_e49fcd23[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ff058abb (
    .a(al_d50b6ef8),
    .b(al_42381c95[7]),
    .c(al_b091d0de[15]),
    .o(al_e49fcd23[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_67444a14 (
    .a(al_d50b6ef8),
    .b(al_42381c95[8]),
    .c(al_b091d0de[16]),
    .o(al_e49fcd23[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a93ef6fc (
    .a(al_d50b6ef8),
    .b(al_42381c95[9]),
    .c(al_b091d0de[17]),
    .o(al_e49fcd23[9]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_d851f814 (
    .a(al_583c216b[0]),
    .b(al_583c216b[3]),
    .c(al_583c216b[5]),
    .d(al_b091d0de[0]),
    .e(al_b091d0de[3]),
    .f(al_b091d0de[5]),
    .o(al_d9d7cf90));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_6b1965f7 (
    .a(al_583c216b[1]),
    .b(al_583c216b[2]),
    .c(al_583c216b[4]),
    .d(al_b091d0de[1]),
    .e(al_b091d0de[2]),
    .f(al_b091d0de[4]),
    .o(al_13db00fa));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    al_3c27dddb (
    .a(al_d9d7cf90),
    .b(al_13db00fa),
    .c(al_583c216b[6]),
    .d(al_b091d0de[6]),
    .o(al_5bd0f2bc));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(~D*~B))"),
    .INIT(32'ha0800a08))
    al_3d8403ac (
    .a(al_5bd0f2bc),
    .b(al_9e8adc84),
    .c(al_583c216b[7]),
    .d(al_96662c62),
    .e(al_b091d0de[7]),
    .o(al_939c27b7));
  AL_DFF_X al_dfd56799 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_939c27b7),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_96662c62));
  AL_MAP_LUT6 #(
    .EQN("(~A*(C*~(B)*~((F*E*~D))+C*B*~((F*E*~D))+~(C)*B*(F*E*~D)+C*B*(F*E*~D)))"),
    .INIT(64'h5044505050505050))
    al_94af0dab (
    .a(al_9e8adc84),
    .b(al_96662c62),
    .c(al_484c4f9e),
    .d(al_7f29f8c[0]),
    .e(al_7f29f8c[1]),
    .f(al_7f29f8c[2]),
    .o(al_feb6df53));
  AL_DFF_X al_25ae3fbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_feb6df53),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_484c4f9e));
  AL_DFF_X al_ec7cd172 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ccdce37d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3910e3c));
  AL_MAP_LUT5 #(
    .EQN("(~D*(E*~(C)*~((B*A))+E*C*~((B*A))+~(E)*C*(B*A)+E*C*(B*A)))"),
    .INIT(32'h00f70080))
    al_b81e6fca (
    .a(al_6f75ef0e),
    .b(rx_clk_en),
    .c(al_4ebb1964),
    .d(al_fea77e50),
    .e(al_a3910e3c),
    .o(al_ccdce37d));
  AL_DFF_0 al_b437afc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[34]));
  AL_DFF_0 al_e9e01220 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[35]));
  AL_DFF_0 al_633a854f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[36]));
  AL_DFF_0 al_8aa99822 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[37]));
  AL_DFF_0 al_4f70c02b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[38]));
  AL_DFF_0 al_b94871 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[39]));
  AL_DFF_0 al_69b5f931 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[40]));
  AL_DFF_0 al_73718271 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[41]));
  AL_DFF_0 al_981c3951 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[42]));
  AL_DFF_0 al_ec608b61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[43]));
  AL_DFF_0 al_76123dff (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[44]));
  AL_DFF_0 al_9b601ad0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[45]));
  AL_DFF_0 al_22d0accb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[46]));
  AL_DFF_0 al_75cde638 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[47]));
  AL_DFF_0 al_4bb3dd9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[48]));
  AL_DFF_0 al_78cffeac (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[49]));
  AL_DFF_0 al_f17caa5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[50]));
  AL_DFF_0 al_3eb413aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[51]));
  AL_DFF_0 al_e0b744f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[52]));
  AL_DFF_0 al_16615310 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[53]));
  AL_DFF_0 al_d73cbbc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[54]));
  AL_DFF_0 al_484cbf68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[55]));
  AL_DFF_0 al_da54a1e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[56]));
  AL_DFF_0 al_f0097b91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[57]));
  AL_DFF_0 al_856b2a0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[58]));
  AL_DFF_0 al_f99e423 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[59]));
  AL_DFF_0 al_8bd52fc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[60]));
  AL_DFF_0 al_9fdf8d1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[61]));
  AL_DFF_0 al_c28e5e67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[62]));
  AL_DFF_0 al_23421334 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[63]));
  AL_DFF_0 al_38bea240 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[0]));
  AL_DFF_0 al_5939186 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[1]));
  AL_DFF_0 al_c8f6d3cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[2]));
  AL_DFF_0 al_7aa32272 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[3]));
  AL_DFF_0 al_718b52e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[4]));
  AL_DFF_0 al_fabf7a6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[5]));
  AL_DFF_0 al_ead28196 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[6]));
  AL_DFF_0 al_ef1a4068 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[7]));
  AL_DFF_0 al_667cf9e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[8]));
  AL_DFF_0 al_ce731eee (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[9]));
  AL_DFF_0 al_80a682a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[10]));
  AL_DFF_0 al_2e06d4bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[11]));
  AL_DFF_0 al_2022ac80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[12]));
  AL_DFF_0 al_93454f14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[13]));
  AL_DFF_0 al_822efda5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[14]));
  AL_DFF_0 al_188edc1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[15]));
  AL_DFF_0 al_eaac19f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[16]));
  AL_DFF_0 al_927f8254 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[17]));
  AL_DFF_0 al_62565de (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[18]));
  AL_DFF_0 al_9bee7d3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[19]));
  AL_DFF_0 al_e786cf59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[20]));
  AL_DFF_0 al_d6dae69e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[21]));
  AL_DFF_0 al_632f271c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[22]));
  AL_DFF_0 al_87838d7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[23]));
  AL_DFF_0 al_1f535962 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[24]));
  AL_DFF_0 al_9987664b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[25]));
  AL_DFF_0 al_7e16e3bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[26]));
  AL_DFF_0 al_af33f630 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[27]));
  AL_DFF_0 al_f2416b3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[28]));
  AL_DFF_0 al_a466055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[29]));
  AL_DFF_0 al_9172742d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[30]));
  AL_DFF_0 al_c8b46f91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_5a460c8d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[31]));
  AL_DFF_0 al_4a06b4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[32]));
  AL_DFF_0 al_dc6a6fe9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_9e004fa1),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_5ffd8cb3[33]));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*D*~C*~B*~A)"),
    .INIT(64'h0000000001000000))
    al_c556b14d (
    .a(s_axi_awaddr[5]),
    .b(s_axi_awaddr[4]),
    .c(s_axi_awaddr[3]),
    .d(s_axi_awaddr[2]),
    .e(s_axi_awaddr[1]),
    .f(s_axi_awaddr[0]),
    .o(al_a9c2861c));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*B*A)"),
    .INIT(32'h08000000))
    al_8fb6fbbc (
    .a(al_a9c2861c),
    .b(s_axi_awaddr[7]),
    .c(s_axi_awaddr[6]),
    .d(s_axi_awvalid),
    .e(s_axi_wvalid),
    .o(al_74d19130));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_68ee2f56 (
    .a(al_74d19130),
    .b(s_axi_wdata[18]),
    .c(al_16296d60),
    .d(al_f931229[2]),
    .o(al_dcfb58ce));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_8e3c87b9 (
    .a(al_74d19130),
    .b(s_axi_wdata[17]),
    .c(al_16296d60),
    .d(al_f931229[1]),
    .o(al_5f4286cf));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_d56e0825 (
    .a(al_74d19130),
    .b(s_axi_wdata[16]),
    .c(al_16296d60),
    .d(al_f931229[0]),
    .o(al_ca35642e));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_586f5bf (
    .a(al_74d19130),
    .b(s_axi_wdata[19]),
    .c(al_16296d60),
    .d(al_f931229[3]),
    .o(al_4276a847));
  AL_DFF_0 al_12c9377c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ca35642e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f931229[0]));
  AL_DFF_0 al_870365d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_5f4286cf),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f931229[1]));
  AL_DFF_0 al_24bf5266 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dcfb58ce),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f931229[2]));
  AL_DFF_0 al_a022cc20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_4276a847),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f931229[3]));
  AL_DFF_X al_1fc5078e (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_593a2319));
  AL_DFF_X al_2740dba9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8dea866b));
  AL_DFF_X al_a8f77686 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f5169e61));
  AL_DFF_X al_b3c0c6f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ee3af5c0));
  AL_DFF_X al_cdeba31d (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_928a2d4f));
  AL_DFF_X al_d935d32f (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5995850b));
  AL_DFF_X al_e670b9a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_70bede4a));
  AL_DFF_X al_bdc98edc (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_58cfbf60));
  AL_DFF_X al_a7a66928 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fe6f17e2));
  AL_DFF_X al_7bf42b6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11243436));
  AL_DFF_X al_25c43df7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b7c18d6c));
  AL_DFF_X al_51c1f1fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f383744d));
  AL_DFF_X al_5c68b4a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8dce46fa));
  AL_DFF_X al_976d69b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_85cd42a7));
  AL_DFF_X al_5c6c8e3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3e863ba));
  AL_DFF_X al_b95a8b87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c55a3d3));
  AL_DFF_X al_68802f91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4cf91e2));
  AL_DFF_X al_1ba3ff11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5d5dee64));
  AL_DFF_X al_101f5a08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7ff105dd));
  AL_DFF_X al_ab3fff10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c32e7d0));
  AL_DFF_X al_2f075d43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e6a1e4d5));
  AL_DFF_X al_b7fd8cd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e2546db0));
  AL_DFF_X al_e1ef64e (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33bf9b84));
  AL_DFF_X al_1babd104 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa8be9ce));
  AL_DFF_X al_412c8dd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f180be0));
  AL_DFF_X al_e8db9cde (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7c64c6fa));
  AL_DFF_X al_94a87418 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe8108));
  AL_DFF_X al_bc760aa0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd2ca50c));
  AL_DFF_X al_6f921b8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b28e21a8));
  AL_DFF_X al_40dc52dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2379dade));
  AL_DFF_X al_ccce065a (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13b54967));
  AL_DFF_X al_37cc0abd (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_b42a6639),
    .d(al_4248a527[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0b71806));
  AL_DFF_X al_299b6c2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_abfa408b[0]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7f29f8c[0]));
  AL_DFF_X al_4c399065 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_abfa408b[1]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7f29f8c[1]));
  AL_DFF_X al_70815a63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_abfa408b[2]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_7f29f8c[2]));
  AL_DFF_X al_8e82abdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[8]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[8]));
  AL_DFF_X al_e1e6ecaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[9]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[9]));
  AL_DFF_X al_63cd5d97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[10]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[10]));
  AL_DFF_X al_c046775b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[11]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[11]));
  AL_DFF_X al_1f49195 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[12]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[12]));
  AL_DFF_X al_fd07ab88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[13]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[13]));
  AL_DFF_X al_6053ac8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[14]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[14]));
  AL_DFF_X al_83d098e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[15]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[15]));
  AL_DFF_X al_34365570 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[16]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[16]));
  AL_DFF_X al_ad026ba2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[17]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[17]));
  AL_DFF_X al_a7b8ca4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[0]));
  AL_DFF_X al_aa3d0960 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[18]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[18]));
  AL_DFF_X al_9054c84b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[19]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[19]));
  AL_DFF_X al_2943f90f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[20]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[20]));
  AL_DFF_X al_b54f968d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[21]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[21]));
  AL_DFF_X al_85aaedef (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[22]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[22]));
  AL_DFF_X al_ad27724 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[23]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[23]));
  AL_DFF_X al_74cadcbc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[24]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[24]));
  AL_DFF_X al_b65efa8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[25]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[25]));
  AL_DFF_X al_c01a616f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[26]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[26]));
  AL_DFF_X al_f7b2f246 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[27]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[27]));
  AL_DFF_X al_63807f8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[1]));
  AL_DFF_X al_41e9847b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[28]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[28]));
  AL_DFF_X al_3ea3aff6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[29]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[29]));
  AL_DFF_X al_7f8e5e44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[30]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[30]));
  AL_DFF_X al_93558748 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[31]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[31]));
  AL_DFF_X al_5053fc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[32]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[32]));
  AL_DFF_X al_45a1bd13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[33]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[33]));
  AL_DFF_X al_d0e1ee5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[34]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[34]));
  AL_DFF_X al_299a8334 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[35]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[35]));
  AL_DFF_X al_77cf9a77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[36]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[36]));
  AL_DFF_X al_ee099ce1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[37]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[37]));
  AL_DFF_X al_707543eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[2]));
  AL_DFF_X al_43c78440 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[38]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[38]));
  AL_DFF_X al_ccc6df58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[39]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[39]));
  AL_DFF_X al_566afcea (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[40]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[40]));
  AL_DFF_X al_8707b74b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[41]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[41]));
  AL_DFF_X al_75d79440 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[42]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[42]));
  AL_DFF_X al_525783c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[43]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[43]));
  AL_DFF_X al_61ee5d83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[44]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[44]));
  AL_DFF_X al_63d4a14e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[45]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[45]));
  AL_DFF_X al_9f535eaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[46]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[46]));
  AL_DFF_X al_eabec868 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[47]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[47]));
  AL_DFF_X al_b63d8636 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[3]));
  AL_DFF_X al_1a453827 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[4]));
  AL_DFF_X al_b7697081 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[5]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[5]));
  AL_DFF_X al_2f3481b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[6]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[6]));
  AL_DFF_X al_cdb2e773 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e49fcd23[7]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b091d0de[7]));
  AL_DFF_0 al_d1aa7c62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[0]));
  AL_DFF_0 al_a58503b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[1]));
  AL_DFF_0 al_3b683095 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[2]));
  AL_DFF_0 al_b312bfea (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[3]));
  AL_DFF_0 al_45c95586 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[4]));
  AL_DFF_0 al_883ca9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[5]));
  AL_DFF_0 al_f9ac9c7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[6]));
  AL_DFF_0 al_fb42ee2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[7]));
  AL_DFF_0 al_36e94ea7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[8]));
  AL_DFF_0 al_cbe47736 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[9]));
  AL_DFF_0 al_88a1d3f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[10]));
  AL_DFF_0 al_69b84d30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[11]));
  AL_DFF_0 al_c7a44bc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[12]));
  AL_DFF_0 al_1e7298f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[13]));
  AL_DFF_0 al_3bd5a832 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[14]));
  AL_DFF_0 al_6167a9ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[15]));
  AL_DFF_0 al_95aa1e3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[16]));
  AL_DFF_0 al_e81310d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[17]));
  AL_DFF_0 al_efc35b7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[18]));
  AL_DFF_0 al_2bbf47ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[19]));
  AL_DFF_0 al_2b370250 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[20]));
  AL_DFF_0 al_42d79268 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[21]));
  AL_DFF_0 al_fa11596f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[22]));
  AL_DFF_0 al_a747a45b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[23]));
  AL_DFF_0 al_811deb27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[24]));
  AL_DFF_0 al_7afbd350 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[25]));
  AL_DFF_0 al_83171202 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[26]));
  AL_DFF_0 al_5f72c58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[27]));
  AL_DFF_0 al_3d37a411 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[28]));
  AL_DFF_0 al_63ecdbde (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[29]));
  AL_DFF_0 al_53151e0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[30]));
  AL_DFF_0 al_d2ee3e73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[31]));
  AL_DFF_0 al_afcd966d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[32]));
  AL_DFF_0 al_1f4a33e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[33]));
  AL_DFF_0 al_f0a04047 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[34]));
  AL_DFF_0 al_c02b34d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[35]));
  AL_DFF_0 al_a53778b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[36]));
  AL_DFF_0 al_fd0e3c43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[37]));
  AL_DFF_0 al_904216e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[38]));
  AL_DFF_0 al_a4da805b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[39]));
  AL_DFF_0 al_3a98b959 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[40]));
  AL_DFF_0 al_b9d7245c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[41]));
  AL_DFF_0 al_fda1b638 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[42]));
  AL_DFF_0 al_73dc1679 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[43]));
  AL_DFF_0 al_4bdfaaf6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[44]));
  AL_DFF_0 al_e86c220b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[45]));
  AL_DFF_0 al_f0afb504 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[46]));
  AL_DFF_0 al_c90128a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ddb70824[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9207c009[47]));
  AL_DFF_X al_be09ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[8]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[8]));
  AL_DFF_X al_13c21e9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[9]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[9]));
  AL_DFF_X al_d999bc57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[10]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[10]));
  AL_DFF_X al_988b1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[11]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[11]));
  AL_DFF_X al_98510ad7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[12]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[12]));
  AL_DFF_X al_47a184b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[13]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[13]));
  AL_DFF_X al_a6c64609 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[14]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[14]));
  AL_DFF_X al_30426b4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[15]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[15]));
  AL_DFF_X al_aabeb068 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[16]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[16]));
  AL_DFF_X al_ea126f78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[17]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[17]));
  AL_DFF_X al_fc13baa8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[0]));
  AL_DFF_X al_8ab73677 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[18]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[18]));
  AL_DFF_X al_9bfa7e95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[19]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[19]));
  AL_DFF_X al_66a9b779 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[20]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[20]));
  AL_DFF_X al_9725663b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[21]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[21]));
  AL_DFF_X al_12e2ce7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[22]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[22]));
  AL_DFF_X al_d7f8b071 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[23]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[23]));
  AL_DFF_X al_91057eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[24]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[24]));
  AL_DFF_X al_f7cc4388 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[25]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[25]));
  AL_DFF_X al_6874f9b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[26]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[26]));
  AL_DFF_X al_36782353 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[27]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[27]));
  AL_DFF_X al_e9a3d81f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[1]));
  AL_DFF_X al_53e47203 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[28]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[28]));
  AL_DFF_X al_e4f007f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[29]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[29]));
  AL_DFF_X al_63f5fb30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[30]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[30]));
  AL_DFF_X al_d7b0a440 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[31]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[31]));
  AL_DFF_X al_95952842 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[32]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[32]));
  AL_DFF_X al_d7657cfb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[33]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[33]));
  AL_DFF_X al_1e4a9cef (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[34]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[34]));
  AL_DFF_X al_3ea01e02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[35]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[35]));
  AL_DFF_X al_4d70f4ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[36]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[36]));
  AL_DFF_X al_4a2f860c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[37]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[37]));
  AL_DFF_X al_dc86438 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[2]));
  AL_DFF_X al_f0527df0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[38]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[38]));
  AL_DFF_X al_c2bc92e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[39]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[39]));
  AL_DFF_X al_599c4ede (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[40]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[40]));
  AL_DFF_X al_937bc85a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[41]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[41]));
  AL_DFF_X al_92bb4d83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[42]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[42]));
  AL_DFF_X al_6b0c1926 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[43]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[43]));
  AL_DFF_X al_8519ca36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[44]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[44]));
  AL_DFF_X al_8371fcae (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[45]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[45]));
  AL_DFF_X al_96070f9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[46]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[46]));
  AL_DFF_X al_7a75bd35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[47]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[47]));
  AL_DFF_X al_ff658fbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[3]));
  AL_DFF_X al_cfb89134 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[4]));
  AL_DFF_X al_18c41e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[5]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[5]));
  AL_DFF_X al_dbc97441 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[6]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[6]));
  AL_DFF_X al_415a2d2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c1c7167[7]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1ef691c[7]));
  AL_DFF_0 al_42324444 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[34]));
  AL_DFF_0 al_312bed8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[35]));
  AL_DFF_0 al_e205d539 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[36]));
  AL_DFF_0 al_ec05de9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[37]));
  AL_DFF_0 al_ccfa9777 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[38]));
  AL_DFF_0 al_8e74f152 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[39]));
  AL_DFF_0 al_e5a3a455 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[40]));
  AL_DFF_0 al_a7c47143 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[41]));
  AL_DFF_0 al_f4098471 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[42]));
  AL_DFF_0 al_ec69e4c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[43]));
  AL_DFF_0 al_aeb8ccb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[44]));
  AL_DFF_0 al_8a43ec7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[45]));
  AL_DFF_0 al_29821fd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[46]));
  AL_DFF_0 al_ea3ab478 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[47]));
  AL_DFF_0 al_fa2243e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[48]));
  AL_DFF_0 al_57293b0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[49]));
  AL_DFF_0 al_f0129e90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[50]));
  AL_DFF_0 al_fec9adfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[51]));
  AL_DFF_0 al_f3e1b3c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[52]));
  AL_DFF_0 al_cf6825ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[53]));
  AL_DFF_0 al_63e7eda1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[54]));
  AL_DFF_0 al_5273df41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[55]));
  AL_DFF_0 al_1bfc5707 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[56]));
  AL_DFF_0 al_b6713c57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[57]));
  AL_DFF_0 al_38f00faf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[58]));
  AL_DFF_0 al_c917bc2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[59]));
  AL_DFF_0 al_18d61af3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[60]));
  AL_DFF_0 al_4ccf9c89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[61]));
  AL_DFF_0 al_5852b80b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[62]));
  AL_DFF_0 al_80cf567b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[63]));
  AL_DFF_0 al_f4fb6aff (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[0]));
  AL_DFF_0 al_c9455f07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[1]));
  AL_DFF_0 al_429f160b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[2]));
  AL_DFF_0 al_6412f607 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[3]));
  AL_DFF_0 al_8be769dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[4]));
  AL_DFF_0 al_23716c2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[5]));
  AL_DFF_0 al_1375f099 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[6]));
  AL_DFF_0 al_b5dd08cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[7]));
  AL_DFF_0 al_f15d6b8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[8]));
  AL_DFF_0 al_c5b6a5e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[9]));
  AL_DFF_0 al_f45cd149 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[10]));
  AL_DFF_0 al_878f51ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[11]));
  AL_DFF_0 al_76932a79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[12]));
  AL_DFF_0 al_d2076f17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[13]));
  AL_DFF_0 al_8d7a25db (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[14]));
  AL_DFF_0 al_926d72c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[15]));
  AL_DFF_0 al_36ce3cbc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[16]));
  AL_DFF_0 al_6e541262 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[17]));
  AL_DFF_0 al_d2ac5d5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[18]));
  AL_DFF_0 al_a1f2a4b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[19]));
  AL_DFF_0 al_82e81999 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[20]));
  AL_DFF_0 al_e64eb7cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[21]));
  AL_DFF_0 al_f4be61b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[22]));
  AL_DFF_0 al_c51e3dd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[23]));
  AL_DFF_0 al_bb888377 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[24]));
  AL_DFF_0 al_e7ff0470 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[25]));
  AL_DFF_0 al_2b13c361 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[26]));
  AL_DFF_0 al_1e18f2eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[27]));
  AL_DFF_0 al_1b502d02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[28]));
  AL_DFF_0 al_79b56aad (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[29]));
  AL_DFF_0 al_f59fc5d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[30]));
  AL_DFF_0 al_5736f9ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_297252e3),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[31]));
  AL_DFF_0 al_bc7298bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[32]));
  AL_DFF_0 al_223a0d8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_db3a7a8b),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_b7012aee[33]));
  AL_DFF_0 al_cfb17be1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[34]));
  AL_DFF_0 al_d09cf1e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[35]));
  AL_DFF_0 al_27c99da3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[36]));
  AL_DFF_0 al_196bb79f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[37]));
  AL_DFF_0 al_1538e47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[38]));
  AL_DFF_0 al_70418e3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[39]));
  AL_DFF_0 al_d38b1705 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[40]));
  AL_DFF_0 al_12bb865f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[41]));
  AL_DFF_0 al_741fca7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[42]));
  AL_DFF_0 al_d4a1d3d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[43]));
  AL_DFF_0 al_e61f7831 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[44]));
  AL_DFF_0 al_496ef118 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[45]));
  AL_DFF_0 al_5113605b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[46]));
  AL_DFF_0 al_ea05ce3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[47]));
  AL_DFF_0 al_56d8d7dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[48]));
  AL_DFF_0 al_8e8faab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[49]));
  AL_DFF_0 al_94f6a133 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[50]));
  AL_DFF_0 al_e9ff23e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[51]));
  AL_DFF_0 al_ab0be9d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[52]));
  AL_DFF_0 al_7f0d399f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[53]));
  AL_DFF_0 al_362fd19d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[54]));
  AL_DFF_0 al_b771a21b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[55]));
  AL_DFF_0 al_13bc854b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[56]));
  AL_DFF_0 al_19b10208 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[57]));
  AL_DFF_0 al_f91c9598 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[58]));
  AL_DFF_0 al_f50b2b4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[59]));
  AL_DFF_0 al_c4aec87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[60]));
  AL_DFF_0 al_1f3f9bb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[61]));
  AL_DFF_0 al_d330d1e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[62]));
  AL_DFF_0 al_5fa8b9ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[63]));
  AL_DFF_0 al_a73af78c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[0]));
  AL_DFF_0 al_36201c6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[1]));
  AL_DFF_0 al_90b8185e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[2]));
  AL_DFF_0 al_16a068ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[3]));
  AL_DFF_0 al_35cb843c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[4]));
  AL_DFF_0 al_a558f70f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[5]));
  AL_DFF_0 al_54344164 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[6]));
  AL_DFF_0 al_9ba8262b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[7]));
  AL_DFF_0 al_e6dbda3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[8]));
  AL_DFF_0 al_d121c0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[9]));
  AL_DFF_0 al_15f97b55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[10]));
  AL_DFF_0 al_433eaf84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[11]));
  AL_DFF_0 al_54f27847 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[12]));
  AL_DFF_0 al_c5db5616 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[13]));
  AL_DFF_0 al_683bc2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[14]));
  AL_DFF_0 al_13c65788 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[15]));
  AL_DFF_0 al_5e92e117 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[16]));
  AL_DFF_0 al_f08e0050 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[17]));
  AL_DFF_0 al_7e561ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[18]));
  AL_DFF_0 al_675e946 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[19]));
  AL_DFF_0 al_69a1715a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[20]));
  AL_DFF_0 al_4b32c9c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[21]));
  AL_DFF_0 al_2272d37b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[22]));
  AL_DFF_0 al_899f0619 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[23]));
  AL_DFF_0 al_612fd227 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[24]));
  AL_DFF_0 al_fd17ddf2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[25]));
  AL_DFF_0 al_4459be40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[26]));
  AL_DFF_0 al_a2645921 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[27]));
  AL_DFF_0 al_4c210943 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[28]));
  AL_DFF_0 al_eb85d76c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[29]));
  AL_DFF_0 al_e332116a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[30]));
  AL_DFF_0 al_f02ecc2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_d0f70766),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[31]));
  AL_DFF_0 al_ed9f4df5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[32]));
  AL_DFF_0 al_2844aaa5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_be4e813d),
    .sr(al_16296d60),
    .ss(1'b0),
    .q(al_f07b9ef6[33]));
  AL_DFF_X al_29492f4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6a2b89f7[3]),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(rx_status_vector[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_45252f80 (
    .a(al_d50b6ef8),
    .b(al_5f463be1),
    .o(al_9e8adc84));
  AL_MAP_LUT6 #(
    .EQN("(~C*~B*~(F@D)*~(E@A))"),
    .INIT(64'h0200010000020001))
    al_402f16c4 (
    .a(al_583c216b[0]),
    .b(al_583c216b[2]),
    .c(al_583c216b[3]),
    .d(al_583c216b[7]),
    .e(al_e8711ae2[0]),
    .f(al_e8711ae2[7]),
    .o(al_abdb8956));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~((~E*D*~C))+~(A)*B*~((~E*D*~C))+A*B*~((~E*D*~C))+~(A)*~(B)*(~E*D*~C)+A*~(B)*(~E*D*~C)+~(A)*B*(~E*D*~C))"),
    .INIT(32'heeeee7ee))
    al_148bfafc (
    .a(al_583c216b[1]),
    .b(al_583c216b[6]),
    .c(al_7f29f8c[0]),
    .d(al_7f29f8c[1]),
    .e(al_7f29f8c[2]),
    .o(al_20628f76));
  AL_MAP_LUT6 #(
    .EQN("(~E*~D*~C*B*~(~F*~A))"),
    .INIT(64'h0000000c00000008))
    al_9c904919 (
    .a(al_9e8adc84),
    .b(al_abdb8956),
    .c(al_20628f76),
    .d(al_583c216b[4]),
    .e(al_583c216b[5]),
    .f(al_8213bac0),
    .o(al_2b4ea789));
  AL_DFF_X al_5301657c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2b4ea789),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_8213bac0));
  AL_MAP_LUT3 #(
    .EQN("(~A*~B*~C+A*~B*C)"),
    .INIT(8'b00100001))
    al_ebe0ef2b (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .o(al_e8711ae2[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~B*~C+~A*B*~C)"),
    .INIT(8'b00000110))
    al_25713970 (
    .a(al_7f29f8c[0]),
    .b(al_7f29f8c[1]),
    .c(al_7f29f8c[2]),
    .o(al_e8711ae2[7]));
  AL_MAP_LUT6 #(
    .EQN("(~A*(E*~(F)*~((D*C*~B))+E*F*~((D*C*~B))+~(E)*F*(D*C*~B)+E*F*(D*C*~B)))"),
    .INIT(64'h5555100045550000))
    al_65fa989a (
    .a(al_9e8adc84),
    .b(al_7f29f8c[0]),
    .c(al_7f29f8c[1]),
    .d(al_7f29f8c[2]),
    .e(al_3aba2254),
    .f(al_8213bac0),
    .o(al_51c4207));
  AL_DFF_X al_915240d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_51c4207),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_3aba2254));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_30c46e18 (
    .a(al_855200e6),
    .b(s_axi_wdata[0]),
    .c(unicast_addr[0]),
    .d(al_16296d60),
    .e(al_9207c009[0]),
    .o(al_ddb70824[0]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_1ab8ec3b (
    .a(al_855200e6),
    .b(s_axi_wdata[10]),
    .c(unicast_addr[10]),
    .d(al_16296d60),
    .e(al_9207c009[10]),
    .o(al_ddb70824[10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_50157d5e (
    .a(al_855200e6),
    .b(s_axi_wdata[11]),
    .c(unicast_addr[11]),
    .d(al_16296d60),
    .e(al_9207c009[11]),
    .o(al_ddb70824[11]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_af54282e (
    .a(al_855200e6),
    .b(s_axi_wdata[12]),
    .c(unicast_addr[12]),
    .d(al_16296d60),
    .e(al_9207c009[12]),
    .o(al_ddb70824[12]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_7cb1c0d2 (
    .a(al_855200e6),
    .b(s_axi_wdata[13]),
    .c(unicast_addr[13]),
    .d(al_16296d60),
    .e(al_9207c009[13]),
    .o(al_ddb70824[13]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_1ca08989 (
    .a(al_855200e6),
    .b(s_axi_wdata[14]),
    .c(unicast_addr[14]),
    .d(al_16296d60),
    .e(al_9207c009[14]),
    .o(al_ddb70824[14]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_58953a0d (
    .a(al_855200e6),
    .b(s_axi_wdata[15]),
    .c(unicast_addr[15]),
    .d(al_16296d60),
    .e(al_9207c009[15]),
    .o(al_ddb70824[15]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_83fc7e59 (
    .a(al_855200e6),
    .b(s_axi_wdata[16]),
    .c(unicast_addr[16]),
    .d(al_16296d60),
    .e(al_9207c009[16]),
    .o(al_ddb70824[16]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_f185842b (
    .a(al_855200e6),
    .b(s_axi_wdata[17]),
    .c(unicast_addr[17]),
    .d(al_16296d60),
    .e(al_9207c009[17]),
    .o(al_ddb70824[17]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_71451622 (
    .a(al_855200e6),
    .b(s_axi_wdata[18]),
    .c(unicast_addr[18]),
    .d(al_16296d60),
    .e(al_9207c009[18]),
    .o(al_ddb70824[18]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_c6b04fce (
    .a(al_855200e6),
    .b(s_axi_wdata[19]),
    .c(unicast_addr[19]),
    .d(al_16296d60),
    .e(al_9207c009[19]),
    .o(al_ddb70824[19]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_48b05f0f (
    .a(al_855200e6),
    .b(s_axi_wdata[1]),
    .c(unicast_addr[1]),
    .d(al_16296d60),
    .e(al_9207c009[1]),
    .o(al_ddb70824[1]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_31751df8 (
    .a(al_855200e6),
    .b(s_axi_wdata[20]),
    .c(unicast_addr[20]),
    .d(al_16296d60),
    .e(al_9207c009[20]),
    .o(al_ddb70824[20]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_3bde1b3b (
    .a(al_855200e6),
    .b(s_axi_wdata[21]),
    .c(unicast_addr[21]),
    .d(al_16296d60),
    .e(al_9207c009[21]),
    .o(al_ddb70824[21]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_2bd94f22 (
    .a(al_855200e6),
    .b(s_axi_wdata[22]),
    .c(unicast_addr[22]),
    .d(al_16296d60),
    .e(al_9207c009[22]),
    .o(al_ddb70824[22]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_a3d904bf (
    .a(al_855200e6),
    .b(s_axi_wdata[23]),
    .c(unicast_addr[23]),
    .d(al_16296d60),
    .e(al_9207c009[23]),
    .o(al_ddb70824[23]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_f4aebe2c (
    .a(al_855200e6),
    .b(s_axi_wdata[24]),
    .c(unicast_addr[24]),
    .d(al_16296d60),
    .e(al_9207c009[24]),
    .o(al_ddb70824[24]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_5e318148 (
    .a(al_855200e6),
    .b(s_axi_wdata[25]),
    .c(unicast_addr[25]),
    .d(al_16296d60),
    .e(al_9207c009[25]),
    .o(al_ddb70824[25]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_4352df1f (
    .a(al_855200e6),
    .b(s_axi_wdata[26]),
    .c(unicast_addr[26]),
    .d(al_16296d60),
    .e(al_9207c009[26]),
    .o(al_ddb70824[26]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_99a811fd (
    .a(al_855200e6),
    .b(s_axi_wdata[27]),
    .c(unicast_addr[27]),
    .d(al_16296d60),
    .e(al_9207c009[27]),
    .o(al_ddb70824[27]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_39bbbe63 (
    .a(al_855200e6),
    .b(s_axi_wdata[28]),
    .c(unicast_addr[28]),
    .d(al_16296d60),
    .e(al_9207c009[28]),
    .o(al_ddb70824[28]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_5fa2fa9c (
    .a(al_855200e6),
    .b(s_axi_wdata[29]),
    .c(unicast_addr[29]),
    .d(al_16296d60),
    .e(al_9207c009[29]),
    .o(al_ddb70824[29]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_d831f27 (
    .a(al_855200e6),
    .b(s_axi_wdata[2]),
    .c(unicast_addr[2]),
    .d(al_16296d60),
    .e(al_9207c009[2]),
    .o(al_ddb70824[2]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_f0e165d7 (
    .a(al_26874532),
    .b(al_60c7c349[0]),
    .c(al_60c7c349[1]),
    .d(al_60c7c349[2]),
    .e(al_60c7c349[3]),
    .o(al_9daabc69));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_40512da5 (
    .a(al_9daabc69),
    .b(al_60c7c349[4]),
    .c(al_60c7c349[5]),
    .d(al_60c7c349[6]),
    .e(al_60c7c349[7]),
    .o(al_855200e6));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_a1bda457 (
    .a(al_855200e6),
    .b(s_axi_wdata[30]),
    .c(unicast_addr[30]),
    .d(al_16296d60),
    .e(al_9207c009[30]),
    .o(al_ddb70824[30]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_29eb6fef (
    .a(al_855200e6),
    .b(s_axi_wdata[31]),
    .c(unicast_addr[31]),
    .d(al_16296d60),
    .e(al_9207c009[31]),
    .o(al_ddb70824[31]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_1347bee0 (
    .a(al_1855fcf8),
    .b(s_axi_wdata[0]),
    .c(unicast_addr[32]),
    .d(al_16296d60),
    .e(al_9207c009[32]),
    .o(al_ddb70824[32]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_72457cb3 (
    .a(al_1855fcf8),
    .b(s_axi_wdata[1]),
    .c(unicast_addr[33]),
    .d(al_16296d60),
    .e(al_9207c009[33]),
    .o(al_ddb70824[33]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_d7b14e9b (
    .a(al_1855fcf8),
    .b(s_axi_wdata[2]),
    .c(unicast_addr[34]),
    .d(al_16296d60),
    .e(al_9207c009[34]),
    .o(al_ddb70824[34]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_f2cfd0ad (
    .a(al_1855fcf8),
    .b(s_axi_wdata[3]),
    .c(unicast_addr[35]),
    .d(al_16296d60),
    .e(al_9207c009[35]),
    .o(al_ddb70824[35]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_e7d28a7e (
    .a(al_1855fcf8),
    .b(s_axi_wdata[4]),
    .c(unicast_addr[36]),
    .d(al_16296d60),
    .e(al_9207c009[36]),
    .o(al_ddb70824[36]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_ea935d81 (
    .a(al_1855fcf8),
    .b(s_axi_wdata[5]),
    .c(unicast_addr[37]),
    .d(al_16296d60),
    .e(al_9207c009[37]),
    .o(al_ddb70824[37]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_6985e40c (
    .a(al_1855fcf8),
    .b(s_axi_wdata[6]),
    .c(unicast_addr[38]),
    .d(al_16296d60),
    .e(al_9207c009[38]),
    .o(al_ddb70824[38]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_4bf18b83 (
    .a(al_1855fcf8),
    .b(s_axi_wdata[7]),
    .c(unicast_addr[39]),
    .d(al_16296d60),
    .e(al_9207c009[39]),
    .o(al_ddb70824[39]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_cbef2940 (
    .a(al_855200e6),
    .b(s_axi_wdata[3]),
    .c(unicast_addr[3]),
    .d(al_16296d60),
    .e(al_9207c009[3]),
    .o(al_ddb70824[3]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_1493e0 (
    .a(al_1855fcf8),
    .b(s_axi_wdata[8]),
    .c(unicast_addr[40]),
    .d(al_16296d60),
    .e(al_9207c009[40]),
    .o(al_ddb70824[40]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_da19ea90 (
    .a(al_1855fcf8),
    .b(s_axi_wdata[9]),
    .c(unicast_addr[41]),
    .d(al_16296d60),
    .e(al_9207c009[41]),
    .o(al_ddb70824[41]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_afa5d9c5 (
    .a(al_1855fcf8),
    .b(s_axi_wdata[10]),
    .c(unicast_addr[42]),
    .d(al_16296d60),
    .e(al_9207c009[42]),
    .o(al_ddb70824[42]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_ce917f3f (
    .a(al_1855fcf8),
    .b(s_axi_wdata[11]),
    .c(unicast_addr[43]),
    .d(al_16296d60),
    .e(al_9207c009[43]),
    .o(al_ddb70824[43]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_408915fa (
    .a(al_1855fcf8),
    .b(s_axi_wdata[12]),
    .c(unicast_addr[44]),
    .d(al_16296d60),
    .e(al_9207c009[44]),
    .o(al_ddb70824[44]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_4443f2e (
    .a(al_1855fcf8),
    .b(s_axi_wdata[13]),
    .c(unicast_addr[45]),
    .d(al_16296d60),
    .e(al_9207c009[45]),
    .o(al_ddb70824[45]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    al_99646d69 (
    .a(al_c9ac0c17),
    .b(al_60c7c349[0]),
    .c(al_60c7c349[1]),
    .d(al_60c7c349[2]),
    .e(al_60c7c349[3]),
    .o(al_1855fcf8));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_501554d0 (
    .a(al_1855fcf8),
    .b(s_axi_wdata[14]),
    .c(unicast_addr[46]),
    .d(al_16296d60),
    .e(al_9207c009[46]),
    .o(al_ddb70824[46]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_b2d771ac (
    .a(al_1855fcf8),
    .b(s_axi_wdata[15]),
    .c(unicast_addr[47]),
    .d(al_16296d60),
    .e(al_9207c009[47]),
    .o(al_ddb70824[47]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_bffdeddd (
    .a(al_855200e6),
    .b(s_axi_wdata[4]),
    .c(unicast_addr[4]),
    .d(al_16296d60),
    .e(al_9207c009[4]),
    .o(al_ddb70824[4]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_d8b2fa59 (
    .a(al_855200e6),
    .b(s_axi_wdata[5]),
    .c(unicast_addr[5]),
    .d(al_16296d60),
    .e(al_9207c009[5]),
    .o(al_ddb70824[5]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_8283d0e4 (
    .a(al_855200e6),
    .b(s_axi_wdata[6]),
    .c(unicast_addr[6]),
    .d(al_16296d60),
    .e(al_9207c009[6]),
    .o(al_ddb70824[6]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_4044e80 (
    .a(al_855200e6),
    .b(s_axi_wdata[7]),
    .c(unicast_addr[7]),
    .d(al_16296d60),
    .e(al_9207c009[7]),
    .o(al_ddb70824[7]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_98012b7f (
    .a(al_855200e6),
    .b(s_axi_wdata[8]),
    .c(unicast_addr[8]),
    .d(al_16296d60),
    .e(al_9207c009[8]),
    .o(al_ddb70824[8]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_1ce6b5e9 (
    .a(al_855200e6),
    .b(s_axi_wdata[9]),
    .c(unicast_addr[9]),
    .d(al_16296d60),
    .e(al_9207c009[9]),
    .o(al_ddb70824[9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dbd91f64 (
    .a(al_d50b6ef8),
    .b(al_9207c009[0]),
    .c(al_f1ef691c[8]),
    .o(al_1c1c7167[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_99e5cef6 (
    .a(al_d50b6ef8),
    .b(al_9207c009[10]),
    .c(al_f1ef691c[18]),
    .o(al_1c1c7167[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e2262b0c (
    .a(al_d50b6ef8),
    .b(al_9207c009[11]),
    .c(al_f1ef691c[19]),
    .o(al_1c1c7167[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5587794a (
    .a(al_d50b6ef8),
    .b(al_9207c009[12]),
    .c(al_f1ef691c[20]),
    .o(al_1c1c7167[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_33ae3b6a (
    .a(al_d50b6ef8),
    .b(al_9207c009[13]),
    .c(al_f1ef691c[21]),
    .o(al_1c1c7167[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4df270a9 (
    .a(al_d50b6ef8),
    .b(al_9207c009[14]),
    .c(al_f1ef691c[22]),
    .o(al_1c1c7167[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6e61f4be (
    .a(al_d50b6ef8),
    .b(al_9207c009[15]),
    .c(al_f1ef691c[23]),
    .o(al_1c1c7167[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bd89be9 (
    .a(al_d50b6ef8),
    .b(al_9207c009[16]),
    .c(al_f1ef691c[24]),
    .o(al_1c1c7167[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_19a101c4 (
    .a(al_d50b6ef8),
    .b(al_9207c009[17]),
    .c(al_f1ef691c[25]),
    .o(al_1c1c7167[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_885b1483 (
    .a(al_d50b6ef8),
    .b(al_9207c009[18]),
    .c(al_f1ef691c[26]),
    .o(al_1c1c7167[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5a066d28 (
    .a(al_d50b6ef8),
    .b(al_9207c009[19]),
    .c(al_f1ef691c[27]),
    .o(al_1c1c7167[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9a474656 (
    .a(al_d50b6ef8),
    .b(al_9207c009[1]),
    .c(al_f1ef691c[9]),
    .o(al_1c1c7167[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c4efb247 (
    .a(al_d50b6ef8),
    .b(al_9207c009[20]),
    .c(al_f1ef691c[28]),
    .o(al_1c1c7167[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b845a603 (
    .a(al_d50b6ef8),
    .b(al_9207c009[21]),
    .c(al_f1ef691c[29]),
    .o(al_1c1c7167[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5662ce7e (
    .a(al_d50b6ef8),
    .b(al_9207c009[22]),
    .c(al_f1ef691c[30]),
    .o(al_1c1c7167[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c27dc281 (
    .a(al_d50b6ef8),
    .b(al_9207c009[23]),
    .c(al_f1ef691c[31]),
    .o(al_1c1c7167[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c5e69592 (
    .a(al_d50b6ef8),
    .b(al_9207c009[24]),
    .c(al_f1ef691c[32]),
    .o(al_1c1c7167[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f87b16ff (
    .a(al_d50b6ef8),
    .b(al_9207c009[25]),
    .c(al_f1ef691c[33]),
    .o(al_1c1c7167[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7850db7 (
    .a(al_d50b6ef8),
    .b(al_9207c009[26]),
    .c(al_f1ef691c[34]),
    .o(al_1c1c7167[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_52710b03 (
    .a(al_d50b6ef8),
    .b(al_9207c009[27]),
    .c(al_f1ef691c[35]),
    .o(al_1c1c7167[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3841a0c (
    .a(al_d50b6ef8),
    .b(al_9207c009[28]),
    .c(al_f1ef691c[36]),
    .o(al_1c1c7167[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8e9a1271 (
    .a(al_d50b6ef8),
    .b(al_9207c009[29]),
    .c(al_f1ef691c[37]),
    .o(al_1c1c7167[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b3d10ac5 (
    .a(al_d50b6ef8),
    .b(al_9207c009[2]),
    .c(al_f1ef691c[10]),
    .o(al_1c1c7167[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_46b9b358 (
    .a(al_d50b6ef8),
    .b(al_9207c009[30]),
    .c(al_f1ef691c[38]),
    .o(al_1c1c7167[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_aae76b99 (
    .a(al_d50b6ef8),
    .b(al_9207c009[31]),
    .c(al_f1ef691c[39]),
    .o(al_1c1c7167[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d13c0da0 (
    .a(al_d50b6ef8),
    .b(al_9207c009[32]),
    .c(al_f1ef691c[40]),
    .o(al_1c1c7167[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2258af64 (
    .a(al_d50b6ef8),
    .b(al_9207c009[33]),
    .c(al_f1ef691c[41]),
    .o(al_1c1c7167[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_de791bb1 (
    .a(al_d50b6ef8),
    .b(al_9207c009[34]),
    .c(al_f1ef691c[42]),
    .o(al_1c1c7167[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_93fa1f55 (
    .a(al_d50b6ef8),
    .b(al_9207c009[35]),
    .c(al_f1ef691c[43]),
    .o(al_1c1c7167[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d64111 (
    .a(al_d50b6ef8),
    .b(al_9207c009[36]),
    .c(al_f1ef691c[44]),
    .o(al_1c1c7167[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a9eabff7 (
    .a(al_d50b6ef8),
    .b(al_9207c009[37]),
    .c(al_f1ef691c[45]),
    .o(al_1c1c7167[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6334a0b7 (
    .a(al_d50b6ef8),
    .b(al_9207c009[38]),
    .c(al_f1ef691c[46]),
    .o(al_1c1c7167[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_21d9b8e2 (
    .a(al_d50b6ef8),
    .b(al_9207c009[39]),
    .c(al_f1ef691c[47]),
    .o(al_1c1c7167[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_10ce9cde (
    .a(al_d50b6ef8),
    .b(al_9207c009[3]),
    .c(al_f1ef691c[11]),
    .o(al_1c1c7167[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_fa28f74b (
    .a(al_d50b6ef8),
    .b(al_9207c009[40]),
    .o(al_1c1c7167[40]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6b2cc39c (
    .a(al_d50b6ef8),
    .b(al_9207c009[41]),
    .o(al_1c1c7167[41]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_7920297e (
    .a(al_d50b6ef8),
    .b(al_9207c009[42]),
    .o(al_1c1c7167[42]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_54b51b14 (
    .a(al_d50b6ef8),
    .b(al_9207c009[43]),
    .o(al_1c1c7167[43]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_4cce180d (
    .a(al_d50b6ef8),
    .b(al_9207c009[44]),
    .o(al_1c1c7167[44]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_cfb3aa3 (
    .a(al_d50b6ef8),
    .b(al_9207c009[45]),
    .o(al_1c1c7167[45]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_afcf3923 (
    .a(al_d50b6ef8),
    .b(al_9207c009[46]),
    .o(al_1c1c7167[46]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_bc081431 (
    .a(al_d50b6ef8),
    .b(al_9207c009[47]),
    .o(al_1c1c7167[47]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_929506fc (
    .a(al_d50b6ef8),
    .b(al_9207c009[4]),
    .c(al_f1ef691c[12]),
    .o(al_1c1c7167[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_635d990f (
    .a(al_d50b6ef8),
    .b(al_9207c009[5]),
    .c(al_f1ef691c[13]),
    .o(al_1c1c7167[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f20b2d23 (
    .a(al_d50b6ef8),
    .b(al_9207c009[6]),
    .c(al_f1ef691c[14]),
    .o(al_1c1c7167[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a2d4c274 (
    .a(al_d50b6ef8),
    .b(al_9207c009[7]),
    .c(al_f1ef691c[15]),
    .o(al_1c1c7167[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6f11b452 (
    .a(al_d50b6ef8),
    .b(al_9207c009[8]),
    .c(al_f1ef691c[16]),
    .o(al_1c1c7167[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_144871ff (
    .a(al_d50b6ef8),
    .b(al_9207c009[9]),
    .c(al_f1ef691c[17]),
    .o(al_1c1c7167[9]));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_af0f831d (
    .a(al_583c216b[2]),
    .b(al_583c216b[3]),
    .c(al_583c216b[5]),
    .d(al_f1ef691c[2]),
    .e(al_f1ef691c[3]),
    .f(al_f1ef691c[5]),
    .o(al_63efbaa0));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(E@B)*~(D@A))"),
    .INIT(64'h8040201008040201))
    al_ad780495 (
    .a(al_583c216b[0]),
    .b(al_583c216b[4]),
    .c(al_583c216b[6]),
    .d(al_f1ef691c[0]),
    .e(al_f1ef691c[4]),
    .f(al_f1ef691c[6]),
    .o(al_6e1ce9f));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    al_866b9848 (
    .a(al_63efbaa0),
    .b(al_6e1ce9f),
    .c(al_583c216b[1]),
    .d(al_f1ef691c[1]),
    .o(al_ae77f168));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D@C)*~(~E*~B))"),
    .INIT(32'ha00a8008))
    al_1a0e3e25 (
    .a(al_ae77f168),
    .b(al_9e8adc84),
    .c(al_583c216b[7]),
    .d(al_f1ef691c[7]),
    .e(al_182d4638),
    .o(al_63cbf333));
  AL_DFF_X al_736bb0bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_63cbf333),
    .en(rx_clk_en),
    .sr(al_fea77e50),
    .ss(1'b0),
    .q(al_182d4638));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_f69628ad (
    .a(al_86bf0006),
    .b(al_c0936433),
    .o(mdio_clk));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_3bf16039 (
    .a(al_6bdd801e),
    .b(al_b2b271cb),
    .c(al_b2deb19c),
    .o(al_51616140));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_22a06ce9 (
    .a(al_51616140),
    .b(al_c99d4c23),
    .o(rx_status_vector[23]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_42d50b03 (
    .a(al_4dabd984),
    .b(al_c99d4c23),
    .c(al_1ce99d34),
    .o(rx_status_vector[24]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_eb655ca8 (
    .a(al_5ffd8cb3[32]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[32]),
    .e(al_f07b9ef6[32]),
    .o(al_98c25345));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_eaec4c0a (
    .a(al_58a4ea01),
    .b(al_98c25345),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_8272529a));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_499dec1c (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[0]),
    .e(al_9207c009[32]),
    .o(al_f5f522a1));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_d062b6cf (
    .a(al_5ffd8cb3[0]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[0]),
    .e(al_f07b9ef6[0]),
    .o(al_bd3e169c));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_bd2cccc1 (
    .a(al_29be6517),
    .b(al_8272529a),
    .c(al_f5f522a1),
    .d(al_bd3e169c),
    .e(al_fa4d6e00[0]),
    .f(al_a927014c),
    .o(al_4248a527[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_c6244f52 (
    .a(al_4248a527[0]),
    .b(al_b42a6639),
    .c(al_2c55a3d3),
    .o(s_axi_rdata[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_a28deb06 (
    .a(al_5ffd8cb3[42]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[42]),
    .e(al_f07b9ef6[42]),
    .o(al_2086e64));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_8b6ab525 (
    .a(al_58a4ea01),
    .b(al_2086e64),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_e739923));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_afa07f72 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[10]),
    .e(al_9207c009[42]),
    .o(al_631f19c6));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_20ff6dac (
    .a(al_5ffd8cb3[10]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[10]),
    .e(al_f07b9ef6[10]),
    .o(al_cad879da));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_43ba4360 (
    .a(al_29be6517),
    .b(al_e739923),
    .c(al_631f19c6),
    .d(al_cad879da),
    .e(al_fa4d6e00[10]),
    .f(al_a927014c),
    .o(al_4248a527[10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_2070e160 (
    .a(al_4248a527[10]),
    .b(al_b42a6639),
    .c(al_7c64c6fa),
    .o(s_axi_rdata[10]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_8cfadf4a (
    .a(al_5ffd8cb3[43]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[43]),
    .e(al_f07b9ef6[43]),
    .o(al_67c63555));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_ebc591e1 (
    .a(al_58a4ea01),
    .b(al_67c63555),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_62f30b7f));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_841b2f96 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[11]),
    .e(al_9207c009[43]),
    .o(al_56607029));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_a7b9b49a (
    .a(al_5ffd8cb3[11]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[11]),
    .e(al_f07b9ef6[11]),
    .o(al_f655e852));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_edfae732 (
    .a(al_29be6517),
    .b(al_62f30b7f),
    .c(al_56607029),
    .d(al_f655e852),
    .e(al_fa4d6e00[11]),
    .f(al_a927014c),
    .o(al_4248a527[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_81b1e95 (
    .a(al_4248a527[11]),
    .b(al_b42a6639),
    .c(al_cafe8108),
    .o(s_axi_rdata[11]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_2f0d60ec (
    .a(al_5ffd8cb3[44]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[44]),
    .e(al_f07b9ef6[44]),
    .o(al_b4de44d1));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_e5710d02 (
    .a(al_58a4ea01),
    .b(al_b4de44d1),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_11c347b2));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_69becd79 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[12]),
    .e(al_9207c009[44]),
    .o(al_581760eb));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_2b4acc64 (
    .a(al_5ffd8cb3[12]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[12]),
    .e(al_f07b9ef6[12]),
    .o(al_c00b14c1));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_fb272503 (
    .a(al_29be6517),
    .b(al_11c347b2),
    .c(al_581760eb),
    .d(al_c00b14c1),
    .e(al_fa4d6e00[12]),
    .f(al_a927014c),
    .o(al_4248a527[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_ab4e6428 (
    .a(al_4248a527[12]),
    .b(al_b42a6639),
    .c(al_cd2ca50c),
    .o(s_axi_rdata[12]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_72fc8a6c (
    .a(al_5ffd8cb3[45]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[45]),
    .e(al_f07b9ef6[45]),
    .o(al_8ae11e67));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_cfb60b14 (
    .a(al_58a4ea01),
    .b(al_8ae11e67),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_c4aea171));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_bc3954b7 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[13]),
    .e(al_9207c009[45]),
    .o(al_b6529d32));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_9e8da5c7 (
    .a(al_5ffd8cb3[13]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[13]),
    .e(al_f07b9ef6[13]),
    .o(al_5ea7feee));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_f0bbb802 (
    .a(al_29be6517),
    .b(al_c4aea171),
    .c(al_b6529d32),
    .d(al_5ea7feee),
    .e(al_fa4d6e00[13]),
    .f(al_a927014c),
    .o(al_4248a527[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_a9c5b70d (
    .a(al_4248a527[13]),
    .b(al_b42a6639),
    .c(al_b28e21a8),
    .o(s_axi_rdata[13]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_343aad73 (
    .a(al_5ffd8cb3[46]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[46]),
    .e(al_f07b9ef6[46]),
    .o(al_414fb589));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_179edb8e (
    .a(al_58a4ea01),
    .b(al_414fb589),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_4753a8f9));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_c66330e (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[14]),
    .e(al_9207c009[46]),
    .o(al_53a5d1d8));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_15cfb9cf (
    .a(al_5ffd8cb3[14]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[14]),
    .e(al_f07b9ef6[14]),
    .o(al_8bc3cc10));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_b6207316 (
    .a(al_29be6517),
    .b(al_4753a8f9),
    .c(al_53a5d1d8),
    .d(al_8bc3cc10),
    .e(al_fa4d6e00[14]),
    .f(al_a927014c),
    .o(al_4248a527[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_cd9e0e06 (
    .a(al_4248a527[14]),
    .b(al_b42a6639),
    .c(al_2379dade),
    .o(s_axi_rdata[14]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_4315d4db (
    .a(al_5ffd8cb3[47]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[47]),
    .e(al_f07b9ef6[47]),
    .o(al_12c00371));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_66d15896 (
    .a(al_58a4ea01),
    .b(al_12c00371),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_68f10ad3));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_e655517a (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[15]),
    .e(al_9207c009[47]),
    .o(al_263a3554));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_c843147a (
    .a(al_5ffd8cb3[15]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[15]),
    .e(al_f07b9ef6[15]),
    .o(al_1cb53946));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_2d598bd1 (
    .a(al_29be6517),
    .b(al_68f10ad3),
    .c(al_263a3554),
    .d(al_1cb53946),
    .e(al_fa4d6e00[15]),
    .f(al_a927014c),
    .o(al_4248a527[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_7a0ed582 (
    .a(al_4248a527[15]),
    .b(al_b42a6639),
    .c(al_13b54967),
    .o(s_axi_rdata[15]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_df829419 (
    .a(al_5ffd8cb3[48]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[48]),
    .e(al_f07b9ef6[48]),
    .o(al_12adcf0d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_459efd44 (
    .a(al_58a4ea01),
    .b(al_12adcf0d),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_a1ae1d55));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_8269a935 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[16]),
    .o(al_38bca4e9));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_a6504da0 (
    .a(al_5ffd8cb3[16]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[16]),
    .e(al_f07b9ef6[16]),
    .o(al_9d0e1a05));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_b9e81c48 (
    .a(al_29be6517),
    .b(al_a1ae1d55),
    .c(al_38bca4e9),
    .d(al_9d0e1a05),
    .e(al_fa4d6e00[16]),
    .f(al_a927014c),
    .o(al_4248a527[16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_6cd9cf62 (
    .a(al_4248a527[16]),
    .b(al_b42a6639),
    .c(al_f0b71806),
    .o(s_axi_rdata[16]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_46da3406 (
    .a(al_5ffd8cb3[49]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[49]),
    .e(al_f07b9ef6[49]),
    .o(al_b6be6226));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_80dca8cd (
    .a(al_58a4ea01),
    .b(al_b6be6226),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_c0e589a5));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_57d4ceec (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[17]),
    .o(al_7bcaf633));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_d97cacc7 (
    .a(al_5ffd8cb3[17]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[17]),
    .e(al_f07b9ef6[17]),
    .o(al_fb677f9));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_53e2b155 (
    .a(al_29be6517),
    .b(al_c0e589a5),
    .c(al_7bcaf633),
    .d(al_fb677f9),
    .e(al_fa4d6e00[17]),
    .f(al_a927014c),
    .o(al_4248a527[17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_17737cb (
    .a(al_4248a527[17]),
    .b(al_b42a6639),
    .c(al_593a2319),
    .o(s_axi_rdata[17]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_1ad35487 (
    .a(al_5ffd8cb3[50]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[50]),
    .e(al_f07b9ef6[50]),
    .o(al_cad59eac));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_561053ac (
    .a(al_58a4ea01),
    .b(al_cad59eac),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_f510713e));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_4f4d2f33 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[18]),
    .o(al_ffaac04));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_627bdcd0 (
    .a(al_5ffd8cb3[18]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[18]),
    .e(al_f07b9ef6[18]),
    .o(al_157db10));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_f30fa362 (
    .a(al_29be6517),
    .b(al_f510713e),
    .c(al_ffaac04),
    .d(al_157db10),
    .e(al_fa4d6e00[18]),
    .f(al_a927014c),
    .o(al_4248a527[18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_45787bba (
    .a(al_4248a527[18]),
    .b(al_b42a6639),
    .c(al_8dea866b),
    .o(s_axi_rdata[18]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_ff898250 (
    .a(al_5ffd8cb3[51]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[51]),
    .e(al_f07b9ef6[51]),
    .o(al_f84368bb));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_1bbb3361 (
    .a(al_58a4ea01),
    .b(al_f84368bb),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_c183d3b1));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_f00b4854 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[19]),
    .o(al_44266b04));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_d9fd072 (
    .a(al_5ffd8cb3[19]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[19]),
    .e(al_f07b9ef6[19]),
    .o(al_a57398e0));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_46d7b34a (
    .a(al_29be6517),
    .b(al_c183d3b1),
    .c(al_44266b04),
    .d(al_a57398e0),
    .e(al_fa4d6e00[19]),
    .f(al_a927014c),
    .o(al_4248a527[19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_5b7960bb (
    .a(al_4248a527[19]),
    .b(al_b42a6639),
    .c(al_f5169e61),
    .o(s_axi_rdata[19]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_22ad3ef7 (
    .a(al_5ffd8cb3[33]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[33]),
    .e(al_f07b9ef6[33]),
    .o(al_b0dc2f75));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_7faf1442 (
    .a(al_58a4ea01),
    .b(al_b0dc2f75),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_e06bf58f));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_82b3a317 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[1]),
    .e(al_9207c009[33]),
    .o(al_ab57e6bf));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_bcb80167 (
    .a(al_5ffd8cb3[1]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[1]),
    .e(al_f07b9ef6[1]),
    .o(al_389c7bee));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_5b81724d (
    .a(al_29be6517),
    .b(al_e06bf58f),
    .c(al_ab57e6bf),
    .d(al_389c7bee),
    .e(al_fa4d6e00[1]),
    .f(al_a927014c),
    .o(al_4248a527[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_a97dfddc (
    .a(al_4248a527[1]),
    .b(al_b42a6639),
    .c(al_e4cf91e2),
    .o(s_axi_rdata[1]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_8a842972 (
    .a(al_5ffd8cb3[52]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[52]),
    .e(al_f07b9ef6[52]),
    .o(al_9149a8cc));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_7c95335f (
    .a(al_58a4ea01),
    .b(al_9149a8cc),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_743eaea9));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_f3ac40bc (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[20]),
    .o(al_5d766886));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_5a9c1d9f (
    .a(al_5ffd8cb3[20]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[20]),
    .e(al_f07b9ef6[20]),
    .o(al_502a557a));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_c43d864 (
    .a(al_29be6517),
    .b(al_743eaea9),
    .c(al_5d766886),
    .d(al_502a557a),
    .e(al_fa4d6e00[20]),
    .f(al_a927014c),
    .o(al_4248a527[20]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b31f66ec (
    .a(al_4248a527[20]),
    .b(al_b42a6639),
    .c(al_ee3af5c0),
    .o(s_axi_rdata[20]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_d820701b (
    .a(al_5ffd8cb3[53]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[53]),
    .e(al_f07b9ef6[53]),
    .o(al_f5fab0c0));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_42e2a628 (
    .a(al_58a4ea01),
    .b(al_f5fab0c0),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_39cac231));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_c32f21fe (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[21]),
    .o(al_429251b));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_3dae4db3 (
    .a(al_5ffd8cb3[21]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[21]),
    .e(al_f07b9ef6[21]),
    .o(al_613f9025));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_bfc904e2 (
    .a(al_29be6517),
    .b(al_39cac231),
    .c(al_429251b),
    .d(al_613f9025),
    .e(al_fa4d6e00[21]),
    .f(al_a927014c),
    .o(al_4248a527[21]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_f9b1c000 (
    .a(al_4248a527[21]),
    .b(al_b42a6639),
    .c(al_928a2d4f),
    .o(s_axi_rdata[21]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_fb3650c1 (
    .a(al_5ffd8cb3[54]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[54]),
    .e(al_f07b9ef6[54]),
    .o(al_6b1e934b));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_fb02fe10 (
    .a(al_58a4ea01),
    .b(al_6b1e934b),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_53e610e6));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_28f8ddd6 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[22]),
    .o(al_8f559a59));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_9f59b362 (
    .a(al_5ffd8cb3[22]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[22]),
    .e(al_f07b9ef6[22]),
    .o(al_43f140b9));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_3c21967f (
    .a(al_29be6517),
    .b(al_53e610e6),
    .c(al_8f559a59),
    .d(al_43f140b9),
    .e(al_fa4d6e00[22]),
    .f(al_a927014c),
    .o(al_4248a527[22]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_f1b90870 (
    .a(al_4248a527[22]),
    .b(al_b42a6639),
    .c(al_5995850b),
    .o(s_axi_rdata[22]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_496e27d7 (
    .a(al_5ffd8cb3[55]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[55]),
    .e(al_f07b9ef6[55]),
    .o(al_3bed0c06));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_c1a46816 (
    .a(al_58a4ea01),
    .b(al_3bed0c06),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_a5ba552b));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_822c8ac8 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[23]),
    .o(al_c246767f));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_cf4fb8ab (
    .a(al_5ffd8cb3[23]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[23]),
    .e(al_f07b9ef6[23]),
    .o(al_43bc4712));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_d8803ef9 (
    .a(al_29be6517),
    .b(al_a5ba552b),
    .c(al_c246767f),
    .d(al_43bc4712),
    .e(al_fa4d6e00[23]),
    .f(al_a927014c),
    .o(al_4248a527[23]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_5ef9b44b (
    .a(al_4248a527[23]),
    .b(al_b42a6639),
    .c(al_70bede4a),
    .o(s_axi_rdata[23]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_2fa7aa45 (
    .a(al_5ffd8cb3[56]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[56]),
    .e(al_f07b9ef6[56]),
    .o(al_82b20445));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_e7e7123f (
    .a(al_58a4ea01),
    .b(al_82b20445),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_d2549f15));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_53f90bb2 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[24]),
    .o(al_6b621a04));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_a1fb098c (
    .a(al_5ffd8cb3[24]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[24]),
    .e(al_f07b9ef6[24]),
    .o(al_c7af49f0));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_58390812 (
    .a(al_29be6517),
    .b(al_d2549f15),
    .c(al_6b621a04),
    .d(al_c7af49f0),
    .e(al_fa4d6e00[24]),
    .f(al_a927014c),
    .o(al_4248a527[24]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_37c2e243 (
    .a(al_4248a527[24]),
    .b(al_b42a6639),
    .c(al_58cfbf60),
    .o(s_axi_rdata[24]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_cbcd87d7 (
    .a(al_5ffd8cb3[57]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[57]),
    .e(al_f07b9ef6[57]),
    .o(al_75607bc2));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_5d3be394 (
    .a(al_58a4ea01),
    .b(al_75607bc2),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_9fedaeeb));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_b5fefc9f (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[25]),
    .o(al_5a10d00d));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_fca5036b (
    .a(al_5ffd8cb3[25]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[25]),
    .e(al_f07b9ef6[25]),
    .o(al_bcfe99bb));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_b6a17aa5 (
    .a(al_29be6517),
    .b(al_9fedaeeb),
    .c(al_5a10d00d),
    .d(al_bcfe99bb),
    .e(al_fa4d6e00[25]),
    .f(al_a927014c),
    .o(al_4248a527[25]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_f129954c (
    .a(al_4248a527[25]),
    .b(al_b42a6639),
    .c(al_fe6f17e2),
    .o(s_axi_rdata[25]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_68614cc7 (
    .a(al_5ffd8cb3[58]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[58]),
    .e(al_f07b9ef6[58]),
    .o(al_40609b11));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_dfa8d1ba (
    .a(al_58a4ea01),
    .b(al_40609b11),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_803791d8));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_727ddd57 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[26]),
    .o(al_f1b5d549));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_c2ee73f6 (
    .a(al_5ffd8cb3[26]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[26]),
    .e(al_f07b9ef6[26]),
    .o(al_67528d08));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_6d25ba7c (
    .a(al_29be6517),
    .b(al_803791d8),
    .c(al_f1b5d549),
    .d(al_67528d08),
    .e(al_fa4d6e00[26]),
    .f(al_a927014c),
    .o(al_4248a527[26]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_7db5613f (
    .a(al_4248a527[26]),
    .b(al_b42a6639),
    .c(al_11243436),
    .o(s_axi_rdata[26]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_74d3877c (
    .a(al_5ffd8cb3[59]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[59]),
    .e(al_f07b9ef6[59]),
    .o(al_54d1791f));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_959a2a4b (
    .a(al_58a4ea01),
    .b(al_54d1791f),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_f75db11b));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_39b65a8f (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[27]),
    .o(al_6ce7e86b));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_cb801194 (
    .a(al_5ffd8cb3[27]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[27]),
    .e(al_f07b9ef6[27]),
    .o(al_2e24cdc2));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_995ccf4 (
    .a(al_29be6517),
    .b(al_f75db11b),
    .c(al_6ce7e86b),
    .d(al_2e24cdc2),
    .e(al_fa4d6e00[27]),
    .f(al_a927014c),
    .o(al_4248a527[27]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_164df7a9 (
    .a(al_4248a527[27]),
    .b(al_b42a6639),
    .c(al_b7c18d6c),
    .o(s_axi_rdata[27]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_1c826caa (
    .a(al_5ffd8cb3[60]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[60]),
    .e(al_f07b9ef6[60]),
    .o(al_ce6f4d2));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_6eae8987 (
    .a(al_58a4ea01),
    .b(al_ce6f4d2),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_899c7875));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_e0cf7dc8 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[28]),
    .o(al_f46dd33d));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_8e81b79 (
    .a(al_5ffd8cb3[28]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[28]),
    .e(al_f07b9ef6[28]),
    .o(al_8868df5f));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_d755193f (
    .a(al_29be6517),
    .b(al_899c7875),
    .c(al_f46dd33d),
    .d(al_8868df5f),
    .e(al_fa4d6e00[28]),
    .f(al_a927014c),
    .o(al_4248a527[28]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e715d086 (
    .a(al_4248a527[28]),
    .b(al_b42a6639),
    .c(al_f383744d),
    .o(s_axi_rdata[28]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_39106382 (
    .a(al_5ffd8cb3[61]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[61]),
    .e(al_f07b9ef6[61]),
    .o(al_816cf877));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_ac798d5b (
    .a(al_58a4ea01),
    .b(al_816cf877),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_83bf8364));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_62cec321 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[29]),
    .o(al_9ca6a99d));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_983df568 (
    .a(al_5ffd8cb3[29]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[29]),
    .e(al_f07b9ef6[29]),
    .o(al_a69b9244));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_c6ecbb87 (
    .a(al_29be6517),
    .b(al_83bf8364),
    .c(al_9ca6a99d),
    .d(al_a69b9244),
    .e(al_fa4d6e00[29]),
    .f(al_a927014c),
    .o(al_4248a527[29]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_27b7c425 (
    .a(al_4248a527[29]),
    .b(al_b42a6639),
    .c(al_8dce46fa),
    .o(s_axi_rdata[29]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_da273e87 (
    .a(al_5ffd8cb3[34]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[34]),
    .e(al_f07b9ef6[34]),
    .o(al_1ca59da3));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_304a754e (
    .a(al_58a4ea01),
    .b(al_1ca59da3),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_f951c654));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_24d2b7a0 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[2]),
    .e(al_9207c009[34]),
    .o(al_4cbbfdff));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_8dffbcdf (
    .a(al_5ffd8cb3[2]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[2]),
    .e(al_f07b9ef6[2]),
    .o(al_6c3542a2));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_afefce (
    .a(al_29be6517),
    .b(al_f951c654),
    .c(al_4cbbfdff),
    .d(al_6c3542a2),
    .e(al_fa4d6e00[2]),
    .f(al_a927014c),
    .o(al_4248a527[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_5267485d (
    .a(al_4248a527[2]),
    .b(al_b42a6639),
    .c(al_5d5dee64),
    .o(s_axi_rdata[2]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_418b67b (
    .a(s_axi_araddr[7]),
    .b(s_axi_araddr[6]),
    .c(s_axi_araddr[5]),
    .d(s_axi_araddr[4]),
    .e(s_axi_araddr[3]),
    .f(s_axi_araddr[0]),
    .o(al_58a4ea01));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_28dc6fcf (
    .a(al_29be6517),
    .b(al_66f1c0a9),
    .c(al_25b9d53e),
    .d(al_2dd67b98),
    .e(al_fa4d6e00[30]),
    .f(al_a927014c),
    .o(al_4248a527[30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e371a3c6 (
    .a(al_4248a527[30]),
    .b(al_b42a6639),
    .c(al_85cd42a7),
    .o(s_axi_rdata[30]));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_f59a983f (
    .a(al_58a4ea01),
    .b(al_a927014c),
    .o(al_b42a6639));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(A*~(~C*B)))"),
    .INIT(32'h0000005d))
    al_b9d63643 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_f931229[2]),
    .e(al_f931229[3]),
    .o(al_29be6517));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_1aa83567 (
    .a(al_5ffd8cb3[62]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[62]),
    .e(al_f07b9ef6[62]),
    .o(al_31b957f1));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_70c3887c (
    .a(al_58a4ea01),
    .b(al_31b957f1),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_66f1c0a9));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_3af804e2 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[30]),
    .o(al_25b9d53e));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_f25b8d97 (
    .a(al_5ffd8cb3[30]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[30]),
    .e(al_f07b9ef6[30]),
    .o(al_2dd67b98));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_5e513d82 (
    .a(al_5ffd8cb3[63]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[63]),
    .e(al_f07b9ef6[63]),
    .o(al_bd973c28));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_39c2b9bb (
    .a(al_58a4ea01),
    .b(al_bd973c28),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_df1c692d));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_5cdd11f3 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[31]),
    .o(al_95b2c02e));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_52332ea1 (
    .a(al_5ffd8cb3[31]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[31]),
    .e(al_f07b9ef6[31]),
    .o(al_a9188fac));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~A*~(~D*B)))*~(F)+~E*(~C*~A*~(~D*B))*~(F)+~(~E)*(~C*~A*~(~D*B))*F+~E*(~C*~A*~(~D*B))*F)"),
    .INIT(64'hfafefafeffff0000))
    al_e7c8e561 (
    .a(al_df1c692d),
    .b(al_29be6517),
    .c(al_95b2c02e),
    .d(al_a9188fac),
    .e(al_fa4d6e00[31]),
    .f(al_a927014c),
    .o(al_4248a527[31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_cf33cdef (
    .a(al_4248a527[31]),
    .b(al_b42a6639),
    .c(al_3e863ba),
    .o(s_axi_rdata[31]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_cff4e5fc (
    .a(al_5ffd8cb3[35]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[35]),
    .e(al_f07b9ef6[35]),
    .o(al_e545d06c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_e1ab61d3 (
    .a(al_58a4ea01),
    .b(al_e545d06c),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_9a8f38a1));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_9754ea1a (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[3]),
    .e(al_9207c009[35]),
    .o(al_6300fa05));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_ca8b616b (
    .a(al_5ffd8cb3[3]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[3]),
    .e(al_f07b9ef6[3]),
    .o(al_93727b8b));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_b0495175 (
    .a(al_29be6517),
    .b(al_9a8f38a1),
    .c(al_6300fa05),
    .d(al_93727b8b),
    .e(al_fa4d6e00[3]),
    .f(al_a927014c),
    .o(al_4248a527[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_972c3cd4 (
    .a(al_4248a527[3]),
    .b(al_b42a6639),
    .c(al_7ff105dd),
    .o(s_axi_rdata[3]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_f77b25a3 (
    .a(al_5ffd8cb3[36]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[36]),
    .e(al_f07b9ef6[36]),
    .o(al_58fac850));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_9e9fc47b (
    .a(al_58a4ea01),
    .b(al_58fac850),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_86319e2));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_565ec14d (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[4]),
    .e(al_9207c009[36]),
    .o(al_842395e3));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_e2bf58c3 (
    .a(al_5ffd8cb3[4]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[4]),
    .e(al_f07b9ef6[4]),
    .o(al_732c5a74));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_54c1faa7 (
    .a(al_29be6517),
    .b(al_86319e2),
    .c(al_842395e3),
    .d(al_732c5a74),
    .e(al_fa4d6e00[4]),
    .f(al_a927014c),
    .o(al_4248a527[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_209c2876 (
    .a(al_4248a527[4]),
    .b(al_b42a6639),
    .c(al_c32e7d0),
    .o(s_axi_rdata[4]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_23f128c8 (
    .a(al_5ffd8cb3[37]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[37]),
    .e(al_f07b9ef6[37]),
    .o(al_d0814789));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_39ae3966 (
    .a(al_58a4ea01),
    .b(al_d0814789),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_b7ea58da));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_bc867d6b (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[5]),
    .e(al_9207c009[37]),
    .o(al_69351137));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_651ab8f6 (
    .a(al_5ffd8cb3[5]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[5]),
    .e(al_f07b9ef6[5]),
    .o(al_5686da25));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_b310d412 (
    .a(al_29be6517),
    .b(al_b7ea58da),
    .c(al_69351137),
    .d(al_5686da25),
    .e(al_fa4d6e00[5]),
    .f(al_a927014c),
    .o(al_4248a527[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_9677aadf (
    .a(al_4248a527[5]),
    .b(al_b42a6639),
    .c(al_e6a1e4d5),
    .o(s_axi_rdata[5]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_a4fbb5bd (
    .a(al_5ffd8cb3[38]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[38]),
    .e(al_f07b9ef6[38]),
    .o(al_1f397d18));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_cb98c06a (
    .a(al_58a4ea01),
    .b(al_1f397d18),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_b723aa66));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_8289f0c6 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[6]),
    .e(al_9207c009[38]),
    .o(al_514ce749));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_922b5b04 (
    .a(al_5ffd8cb3[6]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[6]),
    .e(al_f07b9ef6[6]),
    .o(al_b7dabd2c));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_c28cf809 (
    .a(al_29be6517),
    .b(al_b723aa66),
    .c(al_514ce749),
    .d(al_b7dabd2c),
    .e(al_fa4d6e00[6]),
    .f(al_a927014c),
    .o(al_4248a527[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_3342f245 (
    .a(al_4248a527[6]),
    .b(al_b42a6639),
    .c(al_e2546db0),
    .o(s_axi_rdata[6]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_881b06af (
    .a(al_5ffd8cb3[39]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[39]),
    .e(al_f07b9ef6[39]),
    .o(al_f41510c0));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_c4d98a9b (
    .a(al_58a4ea01),
    .b(al_f41510c0),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_ae9f73b7));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_ade0f96f (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[7]),
    .e(al_9207c009[39]),
    .o(al_b04a4f00));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_7998b693 (
    .a(al_5ffd8cb3[7]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[7]),
    .e(al_f07b9ef6[7]),
    .o(al_74fb81be));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_254667cc (
    .a(al_29be6517),
    .b(al_ae9f73b7),
    .c(al_b04a4f00),
    .d(al_74fb81be),
    .e(al_fa4d6e00[7]),
    .f(al_a927014c),
    .o(al_4248a527[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_7e89b42 (
    .a(al_4248a527[7]),
    .b(al_b42a6639),
    .c(al_33bf9b84),
    .o(s_axi_rdata[7]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_57f29641 (
    .a(al_5ffd8cb3[40]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[40]),
    .e(al_f07b9ef6[40]),
    .o(al_aad3b572));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_85ec254f (
    .a(al_58a4ea01),
    .b(al_aad3b572),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_5039df42));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_1a5830da (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[8]),
    .e(al_9207c009[40]),
    .o(al_5530c5c4));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_bb7d4265 (
    .a(al_5ffd8cb3[8]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[8]),
    .e(al_f07b9ef6[8]),
    .o(al_14a7b701));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_183ce1af (
    .a(al_29be6517),
    .b(al_5039df42),
    .c(al_5530c5c4),
    .d(al_14a7b701),
    .e(al_fa4d6e00[8]),
    .f(al_a927014c),
    .o(al_4248a527[8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_2b83a62a (
    .a(al_4248a527[8]),
    .b(al_b42a6639),
    .c(al_aa8be9ce),
    .o(s_axi_rdata[8]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_6796197b (
    .a(al_5ffd8cb3[41]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[41]),
    .e(al_f07b9ef6[41]),
    .o(al_51967b89));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_2614fc6f (
    .a(al_58a4ea01),
    .b(al_51967b89),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_f931229[2]),
    .f(al_f931229[3]),
    .o(al_40ffa4c8));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_3c421a75 (
    .a(al_58a4ea01),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_9207c009[9]),
    .e(al_9207c009[41]),
    .o(al_70e872b4));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hc1cdf1fd))
    al_9986e1b1 (
    .a(al_5ffd8cb3[9]),
    .b(al_f931229[0]),
    .c(al_f931229[1]),
    .d(al_b7012aee[9]),
    .e(al_f07b9ef6[9]),
    .o(al_fe18e71f));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_ceaf3d78 (
    .a(al_29be6517),
    .b(al_40ffa4c8),
    .c(al_70e872b4),
    .d(al_fe18e71f),
    .e(al_fa4d6e00[9]),
    .f(al_a927014c),
    .o(al_4248a527[9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_f213906a (
    .a(al_4248a527[9]),
    .b(al_b42a6639),
    .c(al_9f180be0),
    .o(s_axi_rdata[9]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_c40e4f13 (
    .a(al_b821ca29),
    .o(speed_1000));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f91da26a (
    .a(speed_100),
    .b(al_b821ca29),
    .o(speed_10));

endmodule 

